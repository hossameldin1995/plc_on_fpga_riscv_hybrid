LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- 00 SW         10
-- 04 KEY        04
-- 08 GPIO_IN    18
-- 0C GPIO_OUT   18
-- 10 LEDG       08
-- 14 LEDR       10

ENTITY Input_Output_Peripheral_REG IS
	PORT( 
		clk		: IN STD_LOGIC;
		reset		: IN STD_LOGIC;
		EN			: IN STD_LOGIC;
		
		KEY		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		LEDR		: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		LEDG		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		SW			: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		
		GPIO_OUT	: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
		GPIO_IN	: IN STD_LOGIC_VECTOR(17 DOWNTO 0);
		
		MW			: IN STD_LOGIC;
		Address	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		IN_Data	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUT_Data	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END;

ARCHITECTURE RTL OF Input_Output_Peripheral_REG IS
	
	SIGNAL LEDR_S		: STD_LOGIC_VECTOR(9 DOWNTO 0);
	SIGNAL LEDG_S		: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL GPIO_OUT_S	: STD_LOGIC_VECTOR(17 DOWNTO 0);
	
	BEGIN
	
	LEDR <= LEDR_S;
	LEDG <= LEDG_S;
	GPIO_OUT <= GPIO_OUT_S;
	
	PROCESS(clk, reset, EN, KEY, SW, GPIO_IN, MW, Address, IN_Data)
	BEGIN
		IF reset = '1' THEN
			GPIO_OUT_S   <= (OTHERS => '0');
			LEDR_S       <= (OTHERS => '0');
			LEDG_S       <= (OTHERS => '0');
			OUT_Data     <= (OTHERS => '0');
		ELSE
			IF EN='1' THEN
				IF MW = '1' then
					IF Address = X"0C" THEN
						GPIO_OUT_S <= IN_Data(17 DOWNTO 0);
					ELSIF Address = X"10" THEN
						LEDG_S <= IN_Data(7 DOWNTO 0);
					ELSIF Address = X"14" THEN
						LEDR_S <= IN_Data(9 DOWNTO 0);
					END IF;
				ELSE -- READ
					IF Address = X"00" THEN
						OUT_Data <= "0000000000000000000000" & SW;
					ELSIF Address = X"04" THEN
						OUT_Data <= "0000000000000000000000000000" & KEY;
					ELSIF Address = X"08" THEN
						OUT_Data <= "00000000000000" & GPIO_IN;
					ELSIF Address = X"0C" THEN
						OUT_Data <= "00000000000000" & GPIO_OUT_S;
					ELSIF Address = X"10" THEN
						OUT_Data <= "000000000000000000000000" & LEDG_S;
					ELSIF Address = X"14" THEN
						OUT_Data <= "0000000000000000000000" & LEDR_S;
					END IF;
				END IF;
			END IF;
		END IF;
	END PROCESS;
END RTL;