----------------------------------------------------------------------------
--! @file
--! @copyright  Copyright 2015 GNSS Sensor Ltd. All right reserved.
--! @author     Sergey Khabarov
--! @brief      Galileo Reference E1 codes.
--! @details    This file contains Galileo E1 codes. (total=32)
--!                  E1c - inav codes  [0..total/2-1]
--!                  E1b - pilot codes [total/2..total-1]
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
--library commonlib;
use work.types_common.all;

entity RomPrn_inferred is
  port (
    clk     : in  std_ulogic;
    inAdr   : in  std_logic_vector(12 downto 0);
    outData : out std_logic_vector(31 downto 0)
  );
end;

architecture rtl of RomPrn_inferred is

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(12 downto 0);

begin

  outData <= romdata;
  
  reg : process (clk) begin
    if rising_edge(clk) then addr <= inAdr; end if;
  end process;
  
  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#0000# => romdata <= X"F5D71013";
    when 16#0001# => romdata <= X"0573541B";
    when 16#0002# => romdata <= X"9DBD4FD9";
    when 16#0003# => romdata <= X"E9B20A0D";
    when 16#0004# => romdata <= X"59D144C5";
    when 16#0005# => romdata <= X"4BC79355";
    when 16#0006# => romdata <= X"39D2E758";
    when 16#0007# => romdata <= X"10FB51E4";
    when 16#0008# => romdata <= X"94093A0A";
    when 16#0009# => romdata <= X"19DD79C7";
    when 16#000A# => romdata <= X"0C5A98E5";
    when 16#000B# => romdata <= X"657AA578";
    when 16#000C# => romdata <= X"097777E8";
    when 16#000D# => romdata <= X"6BCC4651";
    when 16#000E# => romdata <= X"CC72F2F9";
    when 16#000F# => romdata <= X"74DC766E";
    when 16#0010# => romdata <= X"07AEA3D0";
    when 16#0011# => romdata <= X"B557EF42";
    when 16#0012# => romdata <= X"FF57E6A5";
    when 16#0013# => romdata <= X"8E805358";
    when 16#0014# => romdata <= X"CE925766";
    when 16#0015# => romdata <= X"9133B18F";
    when 16#0016# => romdata <= X"80FDBDFB";
    when 16#0017# => romdata <= X"38C5524C";
    when 16#0018# => romdata <= X"7FB1DE07";
    when 16#0019# => romdata <= X"98424829";
    when 16#001A# => romdata <= X"90DF58F7";
    when 16#001B# => romdata <= X"2321D920";
    when 16#001C# => romdata <= X"1F8979EA";
    when 16#001D# => romdata <= X"B159B267";
    when 16#001E# => romdata <= X"9C9E95AA";
    when 16#001F# => romdata <= X"6D53456C";
    when 16#0020# => romdata <= X"0DF75C2B";
    when 16#0021# => romdata <= X"4316D1E2";
    when 16#0022# => romdata <= X"30921688";
    when 16#0023# => romdata <= X"2854253A";
    when 16#0024# => romdata <= X"1FA60CA2";
    when 16#0025# => romdata <= X"C94ECE01";
    when 16#0026# => romdata <= X"3E2A8C94";
    when 16#0027# => romdata <= X"3341E7D9";
    when 16#0028# => romdata <= X"E5A8464B";
    when 16#0029# => romdata <= X"3AD407E0";
    when 16#002A# => romdata <= X"AE465C3E";
    when 16#002B# => romdata <= X"3DD1BE60";
    when 16#002C# => romdata <= X"A8C3D50F";
    when 16#002D# => romdata <= X"83153640";
    when 16#002E# => romdata <= X"1E776BE0";
    when 16#002F# => romdata <= X"2A6042FC";
    when 16#0030# => romdata <= X"4A27AF65";
    when 16#0031# => romdata <= X"3F0CFC4D";
    when 16#0032# => romdata <= X"4D013F11";
    when 16#0033# => romdata <= X"5310788D";
    when 16#0034# => romdata <= X"68CAEAD3";
    when 16#0035# => romdata <= X"ECCCC533";
    when 16#0036# => romdata <= X"0587EB3C";
    when 16#0037# => romdata <= X"22A1459F";
    when 16#0038# => romdata <= X"C8E6FCCE";
    when 16#0039# => romdata <= X"9CDE849A";
    when 16#003A# => romdata <= X"5205E70C";
    when 16#003B# => romdata <= X"6D66D125";
    when 16#003C# => romdata <= X"814D698D";
    when 16#003D# => romdata <= X"D0EEBFEA";
    when 16#003E# => romdata <= X"E52CC65C";
    when 16#003F# => romdata <= X"5C84EEDF";
    when 16#0040# => romdata <= X"20737900";
    when 16#0041# => romdata <= X"0E169D31";
    when 16#0042# => romdata <= X"8426516A";
    when 16#0043# => romdata <= X"C5D1C31F";
    when 16#0044# => romdata <= X"2E18A65E";
    when 16#0045# => romdata <= X"07AE6E33";
    when 16#0046# => romdata <= X"FDD724B1";
    when 16#0047# => romdata <= X"3098B3A4";
    when 16#0048# => romdata <= X"44688389";
    when 16#0049# => romdata <= X"EFBBB5EE";
    when 16#004A# => romdata <= X"AB588742";
    when 16#004B# => romdata <= X"BB083B67";
    when 16#004C# => romdata <= X"9D42FB26";
    when 16#004D# => romdata <= X"FF77919E";
    when 16#004E# => romdata <= X"AB21DE03";
    when 16#004F# => romdata <= X"89D99974";
    when 16#0050# => romdata <= X"98F967AE";
    when 16#0051# => romdata <= X"05AF0F4C";
    when 16#0052# => romdata <= X"7E177416";
    when 16#0053# => romdata <= X"E18C4D5E";
    when 16#0054# => romdata <= X"6987ED35";
    when 16#0055# => romdata <= X"90690AD1";
    when 16#0056# => romdata <= X"27D872F1";
    when 16#0057# => romdata <= X"4A8F4903";
    when 16#0058# => romdata <= X"A1232973";
    when 16#0059# => romdata <= X"2A9768F8";
    when 16#005A# => romdata <= X"2F295BEE";
    when 16#005B# => romdata <= X"39187929";
    when 16#005C# => romdata <= X"3E3A97D5";
    when 16#005D# => romdata <= X"1435A7F0";
    when 16#005E# => romdata <= X"3ED7FBE2";
    when 16#005F# => romdata <= X"75F102A8";
    when 16#0060# => romdata <= X"3202DC3D";
    when 16#0061# => romdata <= X"E94AF4C7";
    when 16#0062# => romdata <= X"12E9D006";
    when 16#0063# => romdata <= X"D182693E";
    when 16#0064# => romdata <= X"9632933E";
    when 16#0065# => romdata <= X"6EB77388";
    when 16#0066# => romdata <= X"0CF147B9";
    when 16#0067# => romdata <= X"22E74539";
    when 16#0068# => romdata <= X"E4582F79";
    when 16#0069# => romdata <= X"E39723B4";
    when 16#006A# => romdata <= X"C80E42ED";
    when 16#006B# => romdata <= X"CE4C08A8";
    when 16#006C# => romdata <= X"D02221BA";
    when 16#006D# => romdata <= X"E6D17734";
    when 16#006E# => romdata <= X"817D5B53";
    when 16#006F# => romdata <= X"1C0D3C1A";
    when 16#0070# => romdata <= X"E723911F";
    when 16#0071# => romdata <= X"3FFF6AAC";
    when 16#0072# => romdata <= X"02E97FEA";
    when 16#0073# => romdata <= X"69E376AF";
    when 16#0074# => romdata <= X"4761E645";
    when 16#0075# => romdata <= X"1CA61FDB";
    when 16#0076# => romdata <= X"2F918764";
    when 16#0077# => romdata <= X"2EFCD63A";
    when 16#0078# => romdata <= X"09AAB680";
    when 16#0079# => romdata <= X"770C1593";
    when 16#007A# => romdata <= X"EEDD4FF4";
    when 16#007B# => romdata <= X"293BFFD6";
    when 16#007C# => romdata <= X"DD2C3367";
    when 16#007D# => romdata <= X"E85B14A6";
    when 16#007E# => romdata <= X"54C834B6";
    when 16#007F# => romdata <= X"699421A0";
    when 16#0080# => romdata <= X"96B856A6";
    when 16#0081# => romdata <= X"29F581D1";
    when 16#0082# => romdata <= X"344FEF59";
    when 16#0083# => romdata <= X"7835FE60";
    when 16#0084# => romdata <= X"434625D0";
    when 16#0085# => romdata <= X"77ECF0D9";
    when 16#0086# => romdata <= X"5FBE1155";
    when 16#0087# => romdata <= X"EA043197";
    when 16#0088# => romdata <= X"9E5AFF54";
    when 16#0089# => romdata <= X"4AF591A3";
    when 16#008A# => romdata <= X"32FDAEF9";
    when 16#008B# => romdata <= X"8AB1EDD8";
    when 16#008C# => romdata <= X"47A73F3A";
    when 16#008D# => romdata <= X"F15AAEE7";
    when 16#008E# => romdata <= X"E9A05C9D";
    when 16#008F# => romdata <= X"82C59EC3";
    when 16#0090# => romdata <= X"25EF4CF2";
    when 16#0091# => romdata <= X"64B8ADF2";
    when 16#0092# => romdata <= X"A8E8BA45";
    when 16#0093# => romdata <= X"9354CB4B";
    when 16#0094# => romdata <= X"415CC50B";
    when 16#0095# => romdata <= X"F239ADBC";
    when 16#0096# => romdata <= X"31B3A9C8";
    when 16#0097# => romdata <= X"7B0843CF";
    when 16#0098# => romdata <= X"3B9E6D64";
    when 16#0099# => romdata <= X"6BA43F86";
    when 16#009A# => romdata <= X"6276B053";
    when 16#009B# => romdata <= X"826F3A23";
    when 16#009C# => romdata <= X"34CC5E2E";
    when 16#009D# => romdata <= X"FB9F8F19";
    when 16#009E# => romdata <= X"5B382E75";
    when 16#009F# => romdata <= X"EEA63F58";
    when 16#00A0# => romdata <= X"A06B3F82";
    when 16#00A1# => romdata <= X"A3B5C77C";
    when 16#00A2# => romdata <= X"1800FD94";
    when 16#00A3# => romdata <= X"98F803E5";
    when 16#00A4# => romdata <= X"24435B32";
    when 16#00A5# => romdata <= X"1210BB84";
    when 16#00A6# => romdata <= X"690BED0B";
    when 16#00A7# => romdata <= X"BBE16D36";
    when 16#00A8# => romdata <= X"3B3A9065";
    when 16#00A9# => romdata <= X"6A73720E";
    when 16#00AA# => romdata <= X"27008852";
    when 16#00AB# => romdata <= X"FB7DACC8";
    when 16#00AC# => romdata <= X"284411B1";
    when 16#00AD# => romdata <= X"77728D95";
    when 16#00AE# => romdata <= X"27C56085";
    when 16#00AF# => romdata <= X"9084A395";
    when 16#00B0# => romdata <= X"A6F11A96";
    when 16#00B1# => romdata <= X"AD9DB6B4";
    when 16#00B2# => romdata <= X"3E00642B";
    when 16#00B3# => romdata <= X"000ED12B";
    when 16#00B4# => romdata <= X"FD967868";
    when 16#00B5# => romdata <= X"EAB11085";
    when 16#00B6# => romdata <= X"52CD4FC8";
    when 16#00B7# => romdata <= X"9FBC408A";
    when 16#00B8# => romdata <= X"CE7678C3";
    when 16#00B9# => romdata <= X"81EC91DD";
    when 16#00BA# => romdata <= X"00031912";
    when 16#00BB# => romdata <= X"4EB5D5EF";
    when 16#00BC# => romdata <= X"52C4CAC9";
    when 16#00BD# => romdata <= X"AADEE2FA";
    when 16#00BE# => romdata <= X"045C16CE";
    when 16#00BF# => romdata <= X"492D7F43";
    when 16#00C0# => romdata <= X"743CA779";
    when 16#00C1# => romdata <= X"24C78696";
    when 16#00C2# => romdata <= X"FCBF2F9F";
    when 16#00C3# => romdata <= X"7F36D8E6";
    when 16#00C4# => romdata <= X"23752200";
    when 16#00C5# => romdata <= X"C6FCBBD7";
    when 16#00C6# => romdata <= X"1ABBB687";
    when 16#00C7# => romdata <= X"7F3C5D6E";
    when 16#00C8# => romdata <= X"6740AB03";
    when 16#00C9# => romdata <= X"89458A6B";
    when 16#00CA# => romdata <= X"66440858";
    when 16#00CB# => romdata <= X"B2D38324";
    when 16#00CC# => romdata <= X"4E853646";
    when 16#00CD# => romdata <= X"FE271421";
    when 16#00CE# => romdata <= X"1DEA9E61";
    when 16#00CF# => romdata <= X"96252815";
    when 16#00D0# => romdata <= X"BB704A20";
    when 16#00D1# => romdata <= X"BFE556AC";
    when 16#00D2# => romdata <= X"474F8998";
    when 16#00D3# => romdata <= X"944E0CAB";
    when 16#00D4# => romdata <= X"BBE21A64";
    when 16#00D5# => romdata <= X"00B87BFD";
    when 16#00D6# => romdata <= X"CF937D12";
    when 16#00D7# => romdata <= X"B2821D59";
    when 16#00D8# => romdata <= X"298AF4AD";
    when 16#00D9# => romdata <= X"378F0F42";
    when 16#00DA# => romdata <= X"BD8C4169";
    when 16#00DB# => romdata <= X"3B8D993C";
    when 16#00DC# => romdata <= X"F37C8B47";
    when 16#00DD# => romdata <= X"8F3BB5D3";
    when 16#00DE# => romdata <= X"3AD2A9FA";
    when 16#00DF# => romdata <= X"24AD7B8F";
    when 16#00E0# => romdata <= X"A895FDBC";
    when 16#00E1# => romdata <= X"04964192";
    when 16#00E2# => romdata <= X"F7BA3FF7";
    when 16#00E3# => romdata <= X"4E0E3A43";
    when 16#00E4# => romdata <= X"5B5DFE04";
    when 16#00E5# => romdata <= X"2E3115CA";
    when 16#00E6# => romdata <= X"CF29624C";
    when 16#00E7# => romdata <= X"0645E9C9";
    when 16#00E8# => romdata <= X"17534A2E";
    when 16#00E9# => romdata <= X"BC1F5665";
    when 16#00EA# => romdata <= X"E4E1B1BC";
    when 16#00EB# => romdata <= X"56208DBC";
    when 16#00EC# => romdata <= X"D8A27CCB";
    when 16#00ED# => romdata <= X"6474D5D0";
    when 16#00EE# => romdata <= X"E20CA407";
    when 16#00EF# => romdata <= X"2C960E5A";
    when 16#00F0# => romdata <= X"CE41BDA3";
    when 16#00F1# => romdata <= X"770DF3B6";
    when 16#00F2# => romdata <= X"81F2B318";
    when 16#00F3# => romdata <= X"F6F8E1CB";
    when 16#00F4# => romdata <= X"17C28573";
    when 16#00F5# => romdata <= X"50FB6009";
    when 16#00F6# => romdata <= X"AED665E1";
    when 16#00F7# => romdata <= X"3B2780D7";
    when 16#00F8# => romdata <= X"9217F73F";
    when 16#00F9# => romdata <= X"AC7A8A48";
    when 16#00FA# => romdata <= X"048DB0FB";
    when 16#00FB# => romdata <= X"8A8A5007";
    when 16#00FC# => romdata <= X"CDDC9A7B";
    when 16#00FD# => romdata <= X"2DA8257C";
    when 16#00FE# => romdata <= X"99F1CB60";
    when 16#00FF# => romdata <= X"5A182040";
    when 16#0100# => romdata <= X"E57DE19A";
    when 16#0101# => romdata <= X"3E4A8C12";
    when 16#0102# => romdata <= X"2FCB1DD6";
    when 16#0103# => romdata <= X"584B3D2D";
    when 16#0104# => romdata <= X"AE364D80";
    when 16#0105# => romdata <= X"0F9C5A9E";
    when 16#0106# => romdata <= X"957B38F6";
    when 16#0107# => romdata <= X"24CBD3AC";
    when 16#0108# => romdata <= X"C58FA3ED";
    when 16#0109# => romdata <= X"070B5E44";
    when 16#010A# => romdata <= X"857CCB81";
    when 16#010B# => romdata <= X"3FBC0BB8";
    when 16#010C# => romdata <= X"3B5D157C";
    when 16#010D# => romdata <= X"6C562422";
    when 16#010E# => romdata <= X"E5963CC4";
    when 16#010F# => romdata <= X"DD753C45";
    when 16#0110# => romdata <= X"B0264F8E";
    when 16#0111# => romdata <= X"136A0F17";
    when 16#0112# => romdata <= X"74D77A54";
    when 16#0113# => romdata <= X"3E44D51E";
    when 16#0114# => romdata <= X"F8C6B940";
    when 16#0115# => romdata <= X"8B6E3B5C";
    when 16#0116# => romdata <= X"EE1347A9";
    when 16#0117# => romdata <= X"4F13ECDC";
    when 16#0118# => romdata <= X"94DC7649";
    when 16#0119# => romdata <= X"76E5A50B";
    when 16#011A# => romdata <= X"4CB0AE75";
    when 16#011B# => romdata <= X"57553B47";
    when 16#011C# => romdata <= X"EDFE03EC";
    when 16#011D# => romdata <= X"2CD32EA8";
    when 16#011E# => romdata <= X"D125A341";
    when 16#011F# => romdata <= X"E1EDFC77";
    when 16#0120# => romdata <= X"E75330D6";
    when 16#0121# => romdata <= X"E7B23DC8";
    when 16#0122# => romdata <= X"38EBCE7E";
    when 16#0123# => romdata <= X"5567F5B8";
    when 16#0124# => romdata <= X"C80C3D15";
    when 16#0125# => romdata <= X"E7404B4E";
    when 16#0126# => romdata <= X"10F0BEB0";
    when 16#0127# => romdata <= X"C69626A8";
    when 16#0128# => romdata <= X"14AF9133";
    when 16#0129# => romdata <= X"4199864F";
    when 16#012A# => romdata <= X"C77E0FF5";
    when 16#012B# => romdata <= X"48DC2A6F";
    when 16#012C# => romdata <= X"A6A71C3C";
    when 16#012D# => romdata <= X"0561F2B0";
    when 16#012E# => romdata <= X"85CC05E8";
    when 16#012F# => romdata <= X"512E27B9";
    when 16#0130# => romdata <= X"DBA60B93";
    when 16#0131# => romdata <= X"D114B879";
    when 16#0132# => romdata <= X"35776C8E";
    when 16#0133# => romdata <= X"9A67905C";
    when 16#0134# => romdata <= X"429D48BF";
    when 16#0135# => romdata <= X"3AB1B0A5";
    when 16#0136# => romdata <= X"6FAFBFD5";
    when 16#0137# => romdata <= X"D9C8D8C8";
    when 16#0138# => romdata <= X"A9E5918B";
    when 16#0139# => romdata <= X"FF273CF5";
    when 16#013A# => romdata <= X"E8664FF2";
    when 16#013B# => romdata <= X"B90314BD";
    when 16#013C# => romdata <= X"BFDAD5AB";
    when 16#013D# => romdata <= X"8C22A0E4";
    when 16#013E# => romdata <= X"5C104ECE";
    when 16#013F# => romdata <= X"75EA43FE";
    when 16#0140# => romdata <= X"9BDCE306";
    when 16#0141# => romdata <= X"A5A28AE4";
    when 16#0142# => romdata <= X"64628163";
    when 16#0143# => romdata <= X"D249D805";
    when 16#0144# => romdata <= X"6005F1A9";
    when 16#0145# => romdata <= X"00951808";
    when 16#0146# => romdata <= X"CC8620F8";
    when 16#0147# => romdata <= X"17681534";
    when 16#0148# => romdata <= X"36F74166";
    when 16#0149# => romdata <= X"7A8E271D";
    when 16#014A# => romdata <= X"D986C7A1";
    when 16#014B# => romdata <= X"E5046FCC";
    when 16#014C# => romdata <= X"74C7CEBB";
    when 16#014D# => romdata <= X"F9A1296D";
    when 16#014E# => romdata <= X"6CF0B2FF";
    when 16#014F# => romdata <= X"85BE412D";
    when 16#0150# => romdata <= X"87214BB3";
    when 16#0151# => romdata <= X"68DFF462";
    when 16#0152# => romdata <= X"AD649D73";
    when 16#0153# => romdata <= X"24A11725";
    when 16#0154# => romdata <= X"2311C664";
    when 16#0155# => romdata <= X"D33E4DAF";
    when 16#0156# => romdata <= X"BD830FBC";
    when 16#0157# => romdata <= X"EB6EFBDD";
    when 16#0158# => romdata <= X"7391D4BA";
    when 16#0159# => romdata <= X"DA7A775F";
    when 16#015A# => romdata <= X"D1949D98";
    when 16#015B# => romdata <= X"1F619655";
    when 16#015C# => romdata <= X"DB3C22BA";
    when 16#015D# => romdata <= X"C34E5AE4";
    when 16#015E# => romdata <= X"1222905C";
    when 16#015F# => romdata <= X"0C7E80D6";
    when 16#0160# => romdata <= X"EA28471E";
    when 16#0161# => romdata <= X"C0468756";
    when 16#0162# => romdata <= X"531C09A4";
    when 16#0163# => romdata <= X"71EDBE20";
    when 16#0164# => romdata <= X"0472E78F";
    when 16#0165# => romdata <= X"1701FEE9";
    when 16#0166# => romdata <= X"6E5769A9";
    when 16#0167# => romdata <= X"893C0F11";
    when 16#0168# => romdata <= X"E7906B06";
    when 16#0169# => romdata <= X"4442E06E";
    when 16#016A# => romdata <= X"21ED8B0D";
    when 16#016B# => romdata <= X"70AF2886";
    when 16#016C# => romdata <= X"90C532A2";
    when 16#016D# => romdata <= X"D03B373E";
    when 16#016E# => romdata <= X"1E0085F6";
    when 16#016F# => romdata <= X"2F7AAA65";
    when 16#0170# => romdata <= X"8B569C51";
    when 16#0171# => romdata <= X"84E3DDC4";
    when 16#0172# => romdata <= X"0ECAA88B";
    when 16#0173# => romdata <= X"88711860";
    when 16#0174# => romdata <= X"1691892F";
    when 16#0175# => romdata <= X"9F55E2DE";
    when 16#0176# => romdata <= X"79E49DFF";
    when 16#0177# => romdata <= X"11D434C2";
    when 16#0178# => romdata <= X"BA3AA644";
    when 16#0179# => romdata <= X"7522A7C9";
    when 16#017A# => romdata <= X"9DC215CA";
    when 16#017B# => romdata <= X"D2ED0114";
    when 16#017C# => romdata <= X"ED62CBDA";
    when 16#017D# => romdata <= X"E9D315E4";
    when 16#017E# => romdata <= X"8AE14D20";
    when 16#017F# => romdata <= X"14B7F8E0";
    when 16#0180# => romdata <= X"C0FC4C72";
    when 16#0181# => romdata <= X"A12023BA";
    when 16#0182# => romdata <= X"7093C867";
    when 16#0183# => romdata <= X"75DF3D2F";
    when 16#0184# => romdata <= X"42C7CEDE";
    when 16#0185# => romdata <= X"61687634";
    when 16#0186# => romdata <= X"0BE43013";
    when 16#0187# => romdata <= X"61B9DC9D";
    when 16#0188# => romdata <= X"FF4F1DEC";
    when 16#0189# => romdata <= X"6A62E165";
    when 16#018A# => romdata <= X"927BDE4F";
    when 16#018B# => romdata <= X"809E969A";
    when 16#018C# => romdata <= X"AD085437";
    when 16#018D# => romdata <= X"496BB959";
    when 16#018E# => romdata <= X"04719820";
    when 16#018F# => romdata <= X"F4CA8ABB";
    when 16#0190# => romdata <= X"A0B84C34";
    when 16#0191# => romdata <= X"B06DD7E2";
    when 16#0192# => romdata <= X"68BA10E3";
    when 16#0193# => romdata <= X"86FA7DB9";
    when 16#0194# => romdata <= X"FCFCDAF2";
    when 16#0195# => romdata <= X"B6AFBA46";
    when 16#0196# => romdata <= X"A8A29915";
    when 16#0197# => romdata <= X"3B4E1158";
    when 16#0198# => romdata <= X"2FBA7F28";
    when 16#0199# => romdata <= X"F0A0F9DE";
    when 16#019A# => romdata <= X"41830AB3";
    when 16#019B# => romdata <= X"3335062C";
    when 16#019C# => romdata <= X"57D81DC3";
    when 16#019D# => romdata <= X"61EDFE49";
    when 16#019E# => romdata <= X"1939100F";
    when 16#019F# => romdata <= X"C827F362";
    when 16#01A0# => romdata <= X"73760043";
    when 16#01A1# => romdata <= X"D1C35B74";
    when 16#01A2# => romdata <= X"E36C6C4D";
    when 16#01A3# => romdata <= X"BE1D3078";
    when 16#01A4# => romdata <= X"47D55AC0";
    when 16#01A5# => romdata <= X"7D8B212C";
    when 16#01A6# => romdata <= X"2DBA632A";
    when 16#01A7# => romdata <= X"86AB15BD";
    when 16#01A8# => romdata <= X"0FAFFA43";
    when 16#01A9# => romdata <= X"070644C7";
    when 16#01AA# => romdata <= X"E5062319";
    when 16#01AB# => romdata <= X"5A3796AA";
    when 16#01AC# => romdata <= X"8E8D6E4E";
    when 16#01AD# => romdata <= X"964FA0E4";
    when 16#01AE# => romdata <= X"488A500B";
    when 16#01AF# => romdata <= X"9063FBBF";
    when 16#01B0# => romdata <= X"B1204A0E";
    when 16#01B1# => romdata <= X"33C6CF28";
    when 16#01B2# => romdata <= X"79AC2BA7";
    when 16#01B3# => romdata <= X"C86CAB57";
    when 16#01B4# => romdata <= X"E3E8A497";
    when 16#01B5# => romdata <= X"836194E6";
    when 16#01B6# => romdata <= X"5C5C39B9";
    when 16#01B7# => romdata <= X"50F1AFC3";
    when 16#01B8# => romdata <= X"B58E850A";
    when 16#01B9# => romdata <= X"5EC39F41";
    when 16#01BA# => romdata <= X"90D55351";
    when 16#01BB# => romdata <= X"D16529CD";
    when 16#01BC# => romdata <= X"52B36DF4";
    when 16#01BD# => romdata <= X"A2DC68EE";
    when 16#01BE# => romdata <= X"202BB758";
    when 16#01BF# => romdata <= X"CF19C54B";
    when 16#01C0# => romdata <= X"0E1461D5";
    when 16#01C1# => romdata <= X"47B5D06C";
    when 16#01C2# => romdata <= X"2F9DC09C";
    when 16#01C3# => romdata <= X"2B15458C";
    when 16#01C4# => romdata <= X"3140860E";
    when 16#01C5# => romdata <= X"4C6F3FE4";
    when 16#01C6# => romdata <= X"F417FDFC";
    when 16#01C7# => romdata <= X"EDE00F71";
    when 16#01C8# => romdata <= X"212EE137";
    when 16#01C9# => romdata <= X"E6669E56";
    when 16#01CA# => romdata <= X"9A784547";
    when 16#01CB# => romdata <= X"0CA564F8";
    when 16#01CC# => romdata <= X"5CB47728";
    when 16#01CD# => romdata <= X"08D65D2B";
    when 16#01CE# => romdata <= X"48D409B7";
    when 16#01CF# => romdata <= X"09BD7AC5";
    when 16#01D0# => romdata <= X"F7E28AA8";
    when 16#01D1# => romdata <= X"04CE9DAC";
    when 16#01D2# => romdata <= X"3ABB5A5B";
    when 16#01D3# => romdata <= X"768C6A18";
    when 16#01D4# => romdata <= X"4B5A974E";
    when 16#01D5# => romdata <= X"933F2C17";
    when 16#01D6# => romdata <= X"72FF64AB";
    when 16#01D7# => romdata <= X"26BA2D5A";
    when 16#01D8# => romdata <= X"165744E3";
    when 16#01D9# => romdata <= X"14EFB223";
    when 16#01DA# => romdata <= X"8AC4858A";
    when 16#01DB# => romdata <= X"8B82723D";
    when 16#01DC# => romdata <= X"AE886547";
    when 16#01DD# => romdata <= X"8EAA261F";
    when 16#01DE# => romdata <= X"35DD4D98";
    when 16#01DF# => romdata <= X"A9C07ACB";
    when 16#01E0# => romdata <= X"0B822AFF";
    when 16#01E1# => romdata <= X"1AD3E739";
    when 16#01E2# => romdata <= X"CB214CE7";
    when 16#01E3# => romdata <= X"37196FEF";
    when 16#01E4# => romdata <= X"2DD0B0D4";
    when 16#01E5# => romdata <= X"5BAC4239";
    when 16#01E6# => romdata <= X"35670BCF";
    when 16#01E7# => romdata <= X"71C2EC04";
    when 16#01E8# => romdata <= X"CCB98943";
    when 16#01E9# => romdata <= X"786173C3";
    when 16#01EA# => romdata <= X"09E75A02";
    when 16#01EB# => romdata <= X"BB78A788";
    when 16#01EC# => romdata <= X"A5E6F8A8";
    when 16#01ED# => romdata <= X"F407E57B";
    when 16#01EE# => romdata <= X"8403841A";
    when 16#01EF# => romdata <= X"9E1FCB3A";
    when 16#01F0# => romdata <= X"7AB80D1F";
    when 16#01F1# => romdata <= X"6529770E";
    when 16#01F2# => romdata <= X"52C173E2";
    when 16#01F3# => romdata <= X"C47EDED4";
    when 16#01F4# => romdata <= X"400D5E66";
    when 16#01F5# => romdata <= X"5E325ED8";
    when 16#01F6# => romdata <= X"45C9E8D0";
    when 16#01F7# => romdata <= X"E66FDA16";
    when 16#01F8# => romdata <= X"B17D61ED";
    when 16#01F9# => romdata <= X"BB336F22";
    when 16#01FA# => romdata <= X"688C3F0F";
    when 16#01FB# => romdata <= X"B040A55F";
    when 16#01FC# => romdata <= X"33B65FA9";
    when 16#01FD# => romdata <= X"F3D45F5B";
    when 16#01FE# => romdata <= X"22C445CB";
    when 16#01FF# => romdata <= X"F9DEB220";
    when 16#0200# => romdata <= X"EA959635";
    when 16#0201# => romdata <= X"7B343DFC";
    when 16#0202# => romdata <= X"31D5875C";
    when 16#0203# => romdata <= X"C0E94117";
    when 16#0204# => romdata <= X"A3365147";
    when 16#0205# => romdata <= X"2E476D38";
    when 16#0206# => romdata <= X"92D8112E";
    when 16#0207# => romdata <= X"B6CB6E01";
    when 16#0208# => romdata <= X"51D409C5";
    when 16#0209# => romdata <= X"A514DCDA";
    when 16#020A# => romdata <= X"38A773C5";
    when 16#020B# => romdata <= X"8F18B590";
    when 16#020C# => romdata <= X"EF9017B6";
    when 16#020D# => romdata <= X"EDF0192A";
    when 16#020E# => romdata <= X"B7EB29DD";
    when 16#020F# => romdata <= X"6E1E7E73";
    when 16#0210# => romdata <= X"90C13E9B";
    when 16#0211# => romdata <= X"10209D57";
    when 16#0212# => romdata <= X"75F3B066";
    when 16#0213# => romdata <= X"F7B2DBB7";
    when 16#0214# => romdata <= X"307FB44F";
    when 16#0215# => romdata <= X"726DD2F3";
    when 16#0216# => romdata <= X"68A5FDBE";
    when 16#0217# => romdata <= X"75BA7248";
    when 16#0218# => romdata <= X"762E1EC7";
    when 16#0219# => romdata <= X"E4589DF1";
    when 16#021A# => romdata <= X"A353A16D";
    when 16#021B# => romdata <= X"6B3CAC1C";
    when 16#021C# => romdata <= X"9ACDB898";
    when 16#021D# => romdata <= X"90ED2C4F";
    when 16#021E# => romdata <= X"44AFEFC7";
    when 16#021F# => romdata <= X"63DB51D1";
    when 16#0220# => romdata <= X"02230C37";
    when 16#0221# => romdata <= X"E1ED0943";
    when 16#0222# => romdata <= X"CD6F4176";
    when 16#0223# => romdata <= X"B2F5C191";
    when 16#0224# => romdata <= X"19588911";
    when 16#0225# => romdata <= X"ACF81A7A";
    when 16#0226# => romdata <= X"29320AD5";
    when 16#0227# => romdata <= X"79C1BFAE";
    when 16#0228# => romdata <= X"D1A70DEE";
    when 16#0229# => romdata <= X"1B870371";
    when 16#022A# => romdata <= X"38ADE411";
    when 16#022B# => romdata <= X"E0BB92F5";
    when 16#022C# => romdata <= X"B3148DFA";
    when 16#022D# => romdata <= X"11F2F84C";
    when 16#022E# => romdata <= X"A6C01912";
    when 16#022F# => romdata <= X"4B922837";
    when 16#0230# => romdata <= X"503AA982";
    when 16#0231# => romdata <= X"3A97E443";
    when 16#0232# => romdata <= X"A66378D5";
    when 16#0233# => romdata <= X"CB3130A7";
    when 16#0234# => romdata <= X"EC9B0567";
    when 16#0235# => romdata <= X"0E85D095";
    when 16#0236# => romdata <= X"D5E6F603";
    when 16#0237# => romdata <= X"092C632E";
    when 16#0238# => romdata <= X"51FD9013";
    when 16#0239# => romdata <= X"FE7FB9F0";
    when 16#023A# => romdata <= X"8448FD09";
    when 16#023B# => romdata <= X"F1219A47";
    when 16#023C# => romdata <= X"44CDAF82";
    when 16#023D# => romdata <= X"BF9C6003";
    when 16#023E# => romdata <= X"9C8185C7";
    when 16#023F# => romdata <= X"E9559FCE";
    when 16#0240# => romdata <= X"301C6D3F";
    when 16#0241# => romdata <= X"46A2E514";
    when 16#0242# => romdata <= X"AAD44D38";
    when 16#0243# => romdata <= X"89C8CB4E";
    when 16#0244# => romdata <= X"D7439BF4";
    when 16#0245# => romdata <= X"7019194F";
    when 16#0246# => romdata <= X"26443637";
    when 16#0247# => romdata <= X"70F8BBD0";
    when 16#0248# => romdata <= X"AE92B6F5";
    when 16#0249# => romdata <= X"F43CBBB5";
    when 16#024A# => romdata <= X"03A88523";
    when 16#024B# => romdata <= X"9DA63690";
    when 16#024C# => romdata <= X"3D4C264B";
    when 16#024D# => romdata <= X"3FF09AB7";
    when 16#024E# => romdata <= X"7E3FDBA7";
    when 16#024F# => romdata <= X"EFC63E07";
    when 16#0250# => romdata <= X"92B6D518";
    when 16#0251# => romdata <= X"3759E57D";
    when 16#0252# => romdata <= X"8A694CDB";
    when 16#0253# => romdata <= X"133B4A9E";
    when 16#0254# => romdata <= X"301CEEEB";
    when 16#0255# => romdata <= X"978050AD";
    when 16#0256# => romdata <= X"9A9E4100";
    when 16#0257# => romdata <= X"91AD29E3";
    when 16#0258# => romdata <= X"89829E2F";
    when 16#0259# => romdata <= X"24BE1E3B";
    when 16#025A# => romdata <= X"24F4540C";
    when 16#025B# => romdata <= X"4A6533EB";
    when 16#025C# => romdata <= X"A72E8AD5";
    when 16#025D# => romdata <= X"40BAAE43";
    when 16#025E# => romdata <= X"A0CB82F9";
    when 16#025F# => romdata <= X"71F3A51D";
    when 16#0260# => romdata <= X"D77FE9E1";
    when 16#0261# => romdata <= X"956E2EE7";
    when 16#0262# => romdata <= X"553E050A";
    when 16#0263# => romdata <= X"1D10B995";
    when 16#0264# => romdata <= X"52DDD5B6";
    when 16#0265# => romdata <= X"8F2E2859";
    when 16#0266# => romdata <= X"712835BD";
    when 16#0267# => romdata <= X"2AD6B088";
    when 16#0268# => romdata <= X"81753B48";
    when 16#0269# => romdata <= X"33FB0474";
    when 16#026A# => romdata <= X"0E3364D2";
    when 16#026B# => romdata <= X"CD4921B9";
    when 16#026C# => romdata <= X"39393E7E";
    when 16#026D# => romdata <= X"A91B854F";
    when 16#026E# => romdata <= X"A1E5A8EE";
    when 16#026F# => romdata <= X"79FF0A83";
    when 16#0270# => romdata <= X"F111F784";
    when 16#0271# => romdata <= X"35481D46";
    when 16#0272# => romdata <= X"2E0E1CBC";
    when 16#0273# => romdata <= X"0C921D19";
    when 16#0274# => romdata <= X"0A435A1B";
    when 16#0275# => romdata <= X"A755E4B7";
    when 16#0276# => romdata <= X"021244FC";
    when 16#0277# => romdata <= X"5E3F0630";
    when 16#0278# => romdata <= X"F2A1F439";
    when 16#0279# => romdata <= X"C02AE619";
    when 16#027A# => romdata <= X"393E5624";
    when 16#027B# => romdata <= X"834B05ED";
    when 16#027C# => romdata <= X"7DEDE5F0";
    when 16#027D# => romdata <= X"AFC7A408";
    when 16#027E# => romdata <= X"99424E75";
    when 16#027F# => romdata <= X"D4EE7920";
    when 16#0280# => romdata <= X"90E92279";
    when 16#0281# => romdata <= X"CD4F60D9";
    when 16#0282# => romdata <= X"8F6E8FCB";
    when 16#0283# => romdata <= X"3E9263DB";
    when 16#0284# => romdata <= X"60FAB146";
    when 16#0285# => romdata <= X"A835AAC2";
    when 16#0286# => romdata <= X"E96B3BE3";
    when 16#0287# => romdata <= X"FF071190";
    when 16#0288# => romdata <= X"32DEE052";
    when 16#0289# => romdata <= X"1C731117";
    when 16#028A# => romdata <= X"E90C2943";
    when 16#028B# => romdata <= X"B389DD6B";
    when 16#028C# => romdata <= X"65C5E21C";
    when 16#028D# => romdata <= X"34F86F5A";
    when 16#028E# => romdata <= X"7ADE0407";
    when 16#028F# => romdata <= X"2DFD1479";
    when 16#0290# => romdata <= X"EA36528D";
    when 16#0291# => romdata <= X"340736B0";
    when 16#0292# => romdata <= X"FED4F620";
    when 16#0293# => romdata <= X"7BE9F6CF";
    when 16#0294# => romdata <= X"C971D5EA";
    when 16#0295# => romdata <= X"11781AC2";
    when 16#0296# => romdata <= X"DA25DBEE";
    when 16#0297# => romdata <= X"B6B903EF";
    when 16#0298# => romdata <= X"8BB0AC0C";
    when 16#0299# => romdata <= X"D2E29F94";
    when 16#029A# => romdata <= X"B8CB6787";
    when 16#029B# => romdata <= X"4A7B7441";
    when 16#029C# => romdata <= X"045758E0";
    when 16#029D# => romdata <= X"9EA06118";
    when 16#029E# => romdata <= X"1A50E0AB";
    when 16#029F# => romdata <= X"7BCCF801";
    when 16#02A0# => romdata <= X"554E0644";
    when 16#02A1# => romdata <= X"780BC137";
    when 16#02A2# => romdata <= X"436E3FB7";
    when 16#02A3# => romdata <= X"784C1828";
    when 16#02A4# => romdata <= X"56A790D6";
    when 16#02A5# => romdata <= X"943BB53D";
    when 16#02A6# => romdata <= X"B40D13D6";
    when 16#02A7# => romdata <= X"A2F7B83A";
    when 16#02A8# => romdata <= X"5C521073";
    when 16#02A9# => romdata <= X"883B90FB";
    when 16#02AA# => romdata <= X"8DB1C0F9";
    when 16#02AB# => romdata <= X"54D13294";
    when 16#02AC# => romdata <= X"3C09156A";
    when 16#02AD# => romdata <= X"09984B82";
    when 16#02AE# => romdata <= X"2079FB8F";
    when 16#02AF# => romdata <= X"D09BC07C";
    when 16#02B0# => romdata <= X"1D6336C7";
    when 16#02B1# => romdata <= X"CEAE8CC3";
    when 16#02B2# => romdata <= X"162760B9";
    when 16#02B3# => romdata <= X"838CA6A3";
    when 16#02B4# => romdata <= X"8FD0044F";
    when 16#02B5# => romdata <= X"DF099E41";
    when 16#02B6# => romdata <= X"6D57BF9F";
    when 16#02B7# => romdata <= X"33A55104";
    when 16#02B8# => romdata <= X"3F34EBF9";
    when 16#02B9# => romdata <= X"BAA90901";
    when 16#02BA# => romdata <= X"E62D2D98";
    when 16#02BB# => romdata <= X"1065F977";
    when 16#02BC# => romdata <= X"852072F6";
    when 16#02BD# => romdata <= X"92535DDE";
    when 16#02BE# => romdata <= X"24EE8946";
    when 16#02BF# => romdata <= X"387B4E5B";
    when 16#02C0# => romdata <= X"0FEFEBD7";
    when 16#02C1# => romdata <= X"5552C1FC";
    when 16#02C2# => romdata <= X"325A608A";
    when 16#02C3# => romdata <= X"78079A9A";
    when 16#02C4# => romdata <= X"C864F2F3";
    when 16#02C5# => romdata <= X"0010A330";
    when 16#02C6# => romdata <= X"4CB16A26";
    when 16#02C7# => romdata <= X"AF98D9BF";
    when 16#02C8# => romdata <= X"D3B8D128";
    when 16#02C9# => romdata <= X"541190B2";
    when 16#02CA# => romdata <= X"BBEE275A";
    when 16#02CB# => romdata <= X"6F53B9BC";
    when 16#02CC# => romdata <= X"51083069";
    when 16#02CD# => romdata <= X"85ECBB98";
    when 16#02CE# => romdata <= X"3B56E34F";
    when 16#02CF# => romdata <= X"18B48A12";
    when 16#02D0# => romdata <= X"AEAB8827";
    when 16#02D1# => romdata <= X"1F4F780C";
    when 16#02D2# => romdata <= X"FDFA83E0";
    when 16#02D3# => romdata <= X"5E35C124";
    when 16#02D4# => romdata <= X"64F43505";
    when 16#02D5# => romdata <= X"97CCAE9B";
    when 16#02D6# => romdata <= X"4498F5A5";
    when 16#02D7# => romdata <= X"454DCC32";
    when 16#02D8# => romdata <= X"18D33367";
    when 16#02D9# => romdata <= X"63674934";
    when 16#02DA# => romdata <= X"ADCBCB5E";
    when 16#02DB# => romdata <= X"A52891EB";
    when 16#02DC# => romdata <= X"240C3622";
    when 16#02DD# => romdata <= X"48226DE6";
    when 16#02DE# => romdata <= X"4899BE30";
    when 16#02DF# => romdata <= X"735F6495";
    when 16#02E0# => romdata <= X"E94AA61A";
    when 16#02E1# => romdata <= X"BEF62B80";
    when 16#02E2# => romdata <= X"3C57FDD0";
    when 16#02E3# => romdata <= X"45B724ED";
    when 16#02E4# => romdata <= X"1966B6E7";
    when 16#02E5# => romdata <= X"DFDFCA5B";
    when 16#02E6# => romdata <= X"36F7B0FA";
    when 16#02E7# => romdata <= X"CEDAC62D";
    when 16#02E8# => romdata <= X"E8E10B12";
    when 16#02E9# => romdata <= X"DFC84B1A";
    when 16#02EA# => romdata <= X"9CEB407B";
    when 16#02EB# => romdata <= X"DE63CDB5";
    when 16#02EC# => romdata <= X"208ABBE5";
    when 16#02ED# => romdata <= X"E066AAF2";
    when 16#02EE# => romdata <= X"62187E94";
    when 16#02EF# => romdata <= X"502B1701";
    when 16#02F0# => romdata <= X"B2CC8681";
    when 16#02F1# => romdata <= X"CB616773";
    when 16#02F2# => romdata <= X"DA2B7AF4";
    when 16#02F3# => romdata <= X"9443CFF5";
    when 16#02F4# => romdata <= X"28F45DD7";
    when 16#02F5# => romdata <= X"F2595983";
    when 16#02F6# => romdata <= X"6771908C";
    when 16#02F7# => romdata <= X"2519171C";
    when 16#02F8# => romdata <= X"AED2BCDC";
    when 16#02F9# => romdata <= X"FCEA4630";
    when 16#02FA# => romdata <= X"1E7D99A5";
    when 16#02FB# => romdata <= X"AF719915";
    when 16#02FC# => romdata <= X"5772E92B";
    when 16#02FD# => romdata <= X"AD85F35E";
    when 16#02FE# => romdata <= X"DB656F09";
    when 16#02FF# => romdata <= X"99EE8280";
    when 16#0300# => romdata <= X"A91F5701";
    when 16#0301# => romdata <= X"02961D62";
    when 16#0302# => romdata <= X"CA6CB551";
    when 16#0303# => romdata <= X"44AFCCEA";
    when 16#0304# => romdata <= X"F3910F33";
    when 16#0305# => romdata <= X"36DCB029";
    when 16#0306# => romdata <= X"CDCBA164";
    when 16#0307# => romdata <= X"ADA72732";
    when 16#0308# => romdata <= X"771B6ECD";
    when 16#0309# => romdata <= X"1C58E49F";
    when 16#030A# => romdata <= X"468A2BFD";
    when 16#030B# => romdata <= X"23E1B996";
    when 16#030C# => romdata <= X"DABABBAF";
    when 16#030D# => romdata <= X"5AB3A4C7";
    when 16#030E# => romdata <= X"4926187B";
    when 16#030F# => romdata <= X"5833006F";
    when 16#0310# => romdata <= X"8BEF7F9C";
    when 16#0311# => romdata <= X"D0F05A2A";
    when 16#0312# => romdata <= X"0B9BD907";
    when 16#0313# => romdata <= X"3C4C3976";
    when 16#0314# => romdata <= X"E8660CE7";
    when 16#0315# => romdata <= X"BF81634C";
    when 16#0316# => romdata <= X"F0B31C3D";
    when 16#0317# => romdata <= X"DD806A6A";
    when 16#0318# => romdata <= X"0C15BC55";
    when 16#0319# => romdata <= X"2B83A867";
    when 16#031A# => romdata <= X"89CC675A";
    when 16#031B# => romdata <= X"6D137BE2";
    when 16#031C# => romdata <= X"7BC86DF6";
    when 16#031D# => romdata <= X"8FEC5D26";
    when 16#031E# => romdata <= X"8119EB9E";
    when 16#031F# => romdata <= X"965260FE";
    when 16#0320# => romdata <= X"1F5C56AE";
    when 16#0321# => romdata <= X"F60A8622";
    when 16#0322# => romdata <= X"CDA8C42F";
    when 16#0323# => romdata <= X"24CBA7F5";
    when 16#0324# => romdata <= X"B07A7416";
    when 16#0325# => romdata <= X"91727732";
    when 16#0326# => romdata <= X"3314AFD3";
    when 16#0327# => romdata <= X"ECD10F74";
    when 16#0328# => romdata <= X"BEE7B22D";
    when 16#0329# => romdata <= X"C760EFA7";
    when 16#032A# => romdata <= X"F935FC99";
    when 16#032B# => romdata <= X"63411353";
    when 16#032C# => romdata <= X"782547FA";
    when 16#032D# => romdata <= X"EED32E69";
    when 16#032E# => romdata <= X"A4FB5756";
    when 16#032F# => romdata <= X"C1A73CCD";
    when 16#0330# => romdata <= X"FFEDE50F";
    when 16#0331# => romdata <= X"4B2D9B5D";
    when 16#0332# => romdata <= X"2ED5C59C";
    when 16#0333# => romdata <= X"9A52D80C";
    when 16#0334# => romdata <= X"D27B989B";
    when 16#0335# => romdata <= X"8DAA14C5";
    when 16#0336# => romdata <= X"69E763C0";
    when 16#0337# => romdata <= X"8FD42358";
    when 16#0338# => romdata <= X"CD064B2D";
    when 16#0339# => romdata <= X"E0526607";
    when 16#033A# => romdata <= X"C9536D75";
    when 16#033B# => romdata <= X"E1617EC8";
    when 16#033C# => romdata <= X"0615EF5E";
    when 16#033D# => romdata <= X"E2314FAC";
    when 16#033E# => romdata <= X"29907B61";
    when 16#033F# => romdata <= X"B61F8696";
    when 16#0340# => romdata <= X"CB80B14B";
    when 16#0341# => romdata <= X"3A0148EE";
    when 16#0342# => romdata <= X"BC825C91";
    when 16#0343# => romdata <= X"150A08A2";
    when 16#0344# => romdata <= X"3FC7B38B";
    when 16#0345# => romdata <= X"5982AA02";
    when 16#0346# => romdata <= X"A18BF6E9";
    when 16#0347# => romdata <= X"1B3A1F2E";
    when 16#0348# => romdata <= X"EF360F68";
    when 16#0349# => romdata <= X"2A34AB36";
    when 16#034A# => romdata <= X"CAFCAD55";
    when 16#034B# => romdata <= X"6841073F";
    when 16#034C# => romdata <= X"219910F7";
    when 16#034D# => romdata <= X"BC2F07CE";
    when 16#034E# => romdata <= X"45E98F77";
    when 16#034F# => romdata <= X"F50475DF";
    when 16#0350# => romdata <= X"9EDFE2DC";
    when 16#0351# => romdata <= X"9E3D7280";
    when 16#0352# => romdata <= X"193D61AB";
    when 16#0353# => romdata <= X"5076A148";
    when 16#0354# => romdata <= X"87E9D919";
    when 16#0355# => romdata <= X"3C3B83C5";
    when 16#0356# => romdata <= X"773BDECA";
    when 16#0357# => romdata <= X"067CA1BC";
    when 16#0358# => romdata <= X"3D4561C3";
    when 16#0359# => romdata <= X"A8B4E300";
    when 16#035A# => romdata <= X"72A6269B";
    when 16#035B# => romdata <= X"529760CA";
    when 16#035C# => romdata <= X"1B5FE9D3";
    when 16#035D# => romdata <= X"DB2B5D12";
    when 16#035E# => romdata <= X"02CE8B18";
    when 16#035F# => romdata <= X"E9E2E80F";
    when 16#0360# => romdata <= X"AFF47108";
    when 16#0361# => romdata <= X"168D3C7E";
    when 16#0362# => romdata <= X"B3C940B1";
    when 16#0363# => romdata <= X"A35A1D1B";
    when 16#0364# => romdata <= X"968A5A9D";
    when 16#0365# => romdata <= X"C0686DD8";
    when 16#0366# => romdata <= X"336E498C";
    when 16#0367# => romdata <= X"240F2087";
    when 16#0368# => romdata <= X"1600FF99";
    when 16#0369# => romdata <= X"5B9E3316";
    when 16#036A# => romdata <= X"9DCFCFCB";
    when 16#036B# => romdata <= X"58E75C94";
    when 16#036C# => romdata <= X"D82F843C";
    when 16#036D# => romdata <= X"60A7118F";
    when 16#036E# => romdata <= X"0D7B4006";
    when 16#036F# => romdata <= X"4A8A4176";
    when 16#0370# => romdata <= X"C5158E86";
    when 16#0371# => romdata <= X"AF0BE4C1";
    when 16#0372# => romdata <= X"D5D73D1C";
    when 16#0373# => romdata <= X"051132A8";
    when 16#0374# => romdata <= X"5CC06284";
    when 16#0375# => romdata <= X"86AFD660";
    when 16#0376# => romdata <= X"502A515D";
    when 16#0377# => romdata <= X"6353B674";
    when 16#0378# => romdata <= X"B1D4E617";
    when 16#0379# => romdata <= X"50C13E8A";
    when 16#037A# => romdata <= X"3AD48FE1";
    when 16#037B# => romdata <= X"F89F201C";
    when 16#037C# => romdata <= X"288A8F44";
    when 16#037D# => romdata <= X"3867C2BA";
    when 16#037E# => romdata <= X"C23C706E";
    when 16#037F# => romdata <= X"E7A2D2C0";
    when 16#0380# => romdata <= X"C6E00978";
    when 16#0381# => romdata <= X"E3511645";
    when 16#0382# => romdata <= X"32EEA256";
    when 16#0383# => romdata <= X"ECBE0D4F";
    when 16#0384# => romdata <= X"8FCE02A2";
    when 16#0385# => romdata <= X"76BD1966";
    when 16#0386# => romdata <= X"6DE93936";
    when 16#0387# => romdata <= X"F7A242FC";
    when 16#0388# => romdata <= X"4C7E8797";
    when 16#0389# => romdata <= X"91314B04";
    when 16#038A# => romdata <= X"3ABF1D5F";
    when 16#038B# => romdata <= X"9B0036ED";
    when 16#038C# => romdata <= X"22AA9202";
    when 16#038D# => romdata <= X"8C800C4D";
    when 16#038E# => romdata <= X"62BD6640";
    when 16#038F# => romdata <= X"431170EA";
    when 16#0390# => romdata <= X"77311865";
    when 16#0391# => romdata <= X"074D670A";
    when 16#0392# => romdata <= X"F2847AA4";
    when 16#0393# => romdata <= X"7CB94584";
    when 16#0394# => romdata <= X"A793FA82";
    when 16#0395# => romdata <= X"F51574BD";
    when 16#0396# => romdata <= X"7C62BF14";
    when 16#0397# => romdata <= X"386F14A3";
    when 16#0398# => romdata <= X"D7DBD129";
    when 16#0399# => romdata <= X"FDE64EAD";
    when 16#039A# => romdata <= X"67EB35D5";
    when 16#039B# => romdata <= X"E13FF214";
    when 16#039C# => romdata <= X"D7D163B7";
    when 16#039D# => romdata <= X"70D4A77A";
    when 16#039E# => romdata <= X"62D02D88";
    when 16#039F# => romdata <= X"C0FCF3FA";
    when 16#03A0# => romdata <= X"5EC306EB";
    when 16#03A1# => romdata <= X"7F855391";
    when 16#03A2# => romdata <= X"05FA2CE5";
    when 16#03A3# => romdata <= X"F53D182E";
    when 16#03A4# => romdata <= X"58FBBC1C";
    when 16#03A5# => romdata <= X"57CFBCD2";
    when 16#03A6# => romdata <= X"D2F7FC8A";
    when 16#03A7# => romdata <= X"067D6FA0";
    when 16#03A8# => romdata <= X"BC834DAB";
    when 16#03A9# => romdata <= X"8F370B09";
    when 16#03AA# => romdata <= X"71BF6D06";
    when 16#03AB# => romdata <= X"8CD4D3A3";
    when 16#03AC# => romdata <= X"2C11C659";
    when 16#03AD# => romdata <= X"8DEBBAEA";
    when 16#03AE# => romdata <= X"046528C5";
    when 16#03AF# => romdata <= X"EF762828";
    when 16#03B0# => romdata <= X"CC84D003";
    when 16#03B1# => romdata <= X"847069FA";
    when 16#03B2# => romdata <= X"18743A80";
    when 16#03B3# => romdata <= X"9A004431";
    when 16#03B4# => romdata <= X"E83924B8";
    when 16#03B5# => romdata <= X"FDF0AC78";
    when 16#03B6# => romdata <= X"699B905A";
    when 16#03B7# => romdata <= X"CCFF82E8";
    when 16#03B8# => romdata <= X"3FDAFEC8";
    when 16#03B9# => romdata <= X"648DF640";
    when 16#03BA# => romdata <= X"42FC9438";
    when 16#03BB# => romdata <= X"B261B73F";
    when 16#03BC# => romdata <= X"0541498A";
    when 16#03BD# => romdata <= X"CAD67D70";
    when 16#03BE# => romdata <= X"2AB631BE";
    when 16#03BF# => romdata <= X"CEF8680D";
    when 16#03C0# => romdata <= X"33CE8F4F";
    when 16#03C1# => romdata <= X"0CE29B95";
    when 16#03C2# => romdata <= X"132591A3";
    when 16#03C3# => romdata <= X"50DD68B3";
    when 16#03C4# => romdata <= X"6734B97D";
    when 16#03C5# => romdata <= X"4B3E84A7";
    when 16#03C6# => romdata <= X"6497F702";
    when 16#03C7# => romdata <= X"312F2A83";
    when 16#03C8# => romdata <= X"70DCF26A";
    when 16#03C9# => romdata <= X"7C3C8EB9";
    when 16#03CA# => romdata <= X"1DD8699C";
    when 16#03CB# => romdata <= X"48F55175";
    when 16#03CC# => romdata <= X"0712683E";
    when 16#03CD# => romdata <= X"03970837";
    when 16#03CE# => romdata <= X"14A6CAC3";
    when 16#03CF# => romdata <= X"457C0FA7";
    when 16#03D0# => romdata <= X"0BB3A036";
    when 16#03D1# => romdata <= X"C6E0BEF2";
    when 16#03D2# => romdata <= X"4E6B20BA";
    when 16#03D3# => romdata <= X"5565B351";
    when 16#03D4# => romdata <= X"C2EFD56B";
    when 16#03D5# => romdata <= X"D9455FF7";
    when 16#03D6# => romdata <= X"728BE07A";
    when 16#03D7# => romdata <= X"097208E7";
    when 16#03D8# => romdata <= X"3DE4CD0C";
    when 16#03D9# => romdata <= X"B4E215B4";
    when 16#03DA# => romdata <= X"64236512";
    when 16#03DB# => romdata <= X"3CDEA419";
    when 16#03DC# => romdata <= X"B28459D5";
    when 16#03DD# => romdata <= X"0E864B76";
    when 16#03DE# => romdata <= X"2554E7C1";
    when 16#03DF# => romdata <= X"D7CAF73D";
    when 16#03E0# => romdata <= X"A7D40EDE";
    when 16#03E1# => romdata <= X"F5D824A2";
    when 16#03E2# => romdata <= X"FE1A6CA4";
    when 16#03E3# => romdata <= X"73B07370";
    when 16#03E4# => romdata <= X"932A8A5D";
    when 16#03E5# => romdata <= X"441DEE3C";
    when 16#03E6# => romdata <= X"9A60DB68";
    when 16#03E7# => romdata <= X"E27A9D3E";
    when 16#03E8# => romdata <= X"9C8229B4";
    when 16#03E9# => romdata <= X"4E5B434C";
    when 16#03EA# => romdata <= X"6D18A8CA";
    when 16#03EB# => romdata <= X"DB6D17BC";
    when 16#03EC# => romdata <= X"4614DEBE";
    when 16#03ED# => romdata <= X"AD670C73";
    when 16#03EE# => romdata <= X"132CE2F9";
    when 16#03EF# => romdata <= X"99C8716D";
    when 16#03F0# => romdata <= X"1098C692";
    when 16#03F1# => romdata <= X"77E8ECAC";
    when 16#03F2# => romdata <= X"546EF800";
    when 16#03F3# => romdata <= X"2E5182E2";
    when 16#03F4# => romdata <= X"5F31A354";
    when 16#03F5# => romdata <= X"DF112E97";
    when 16#03F6# => romdata <= X"F8733DD2";
    when 16#03F7# => romdata <= X"0893B430";
    when 16#03F8# => romdata <= X"CD7130E6";
    when 16#03F9# => romdata <= X"9ED4A0FE";
    when 16#03FA# => romdata <= X"4D6C2E4F";
    when 16#03FB# => romdata <= X"A479001E";
    when 16#03FC# => romdata <= X"42EBC9F3";
    when 16#03FD# => romdata <= X"6E5DFD3E";
    when 16#03FE# => romdata <= X"0BE35A64";
    when 16#03FF# => romdata <= X"B89745E0";
    when 16#0400# => romdata <= X"821BBB3F";
    when 16#0401# => romdata <= X"B91E5025";
    when 16#0402# => romdata <= X"3A9E71AC";
    when 16#0403# => romdata <= X"379ED57A";
    when 16#0404# => romdata <= X"EF394C2C";
    when 16#0405# => romdata <= X"C59587B2";
    when 16#0406# => romdata <= X"D0337CE7";
    when 16#0407# => romdata <= X"4002EEAD";
    when 16#0408# => romdata <= X"17AB5D50";
    when 16#0409# => romdata <= X"4BCA68BD";
    when 16#040A# => romdata <= X"AE9061C3";
    when 16#040B# => romdata <= X"DBAE2985";
    when 16#040C# => romdata <= X"EBE292B9";
    when 16#040D# => romdata <= X"BEC9D354";
    when 16#040E# => romdata <= X"2015225F";
    when 16#040F# => romdata <= X"44ED3C2C";
    when 16#0410# => romdata <= X"3FFB036A";
    when 16#0411# => romdata <= X"515BF33D";
    when 16#0412# => romdata <= X"A1690F34";
    when 16#0413# => romdata <= X"38FD225A";
    when 16#0414# => romdata <= X"5034106C";
    when 16#0415# => romdata <= X"5F4BCC43";
    when 16#0416# => romdata <= X"301EEC22";
    when 16#0417# => romdata <= X"45D73F63";
    when 16#0418# => romdata <= X"038E2A7D";
    when 16#0419# => romdata <= X"9B8CF95A";
    when 16#041A# => romdata <= X"9FD813FF";
    when 16#041B# => romdata <= X"A071FFDE";
    when 16#041C# => romdata <= X"423E0CE7";
    when 16#041D# => romdata <= X"37969578";
    when 16#041E# => romdata <= X"BEB90976";
    when 16#041F# => romdata <= X"4A8D6DAA";
    when 16#0420# => romdata <= X"9E15A4FA";
    when 16#0421# => romdata <= X"08678316";
    when 16#0422# => romdata <= X"52C0F6E9";
    when 16#0423# => romdata <= X"AAA39A63";
    when 16#0424# => romdata <= X"F0AEEF62";
    when 16#0425# => romdata <= X"A433476C";
    when 16#0426# => romdata <= X"C7380460";
    when 16#0427# => romdata <= X"ECFB8B7F";
    when 16#0428# => romdata <= X"3B2FE8C4";
    when 16#0429# => romdata <= X"C42A3EF1";
    when 16#042A# => romdata <= X"CDB808FC";
    when 16#042B# => romdata <= X"9747FB4F";
    when 16#042C# => romdata <= X"044B3B47";
    when 16#042D# => romdata <= X"A4EDFCC9";
    when 16#042E# => romdata <= X"463ABB72";
    when 16#042F# => romdata <= X"C55399B2";
    when 16#0430# => romdata <= X"F79EE5FE";
    when 16#0431# => romdata <= X"DA270D63";
    when 16#0432# => romdata <= X"58B27F84";
    when 16#0433# => romdata <= X"66969DE4";
    when 16#0434# => romdata <= X"A5F2E6A5";
    when 16#0435# => romdata <= X"F2C4CF08";
    when 16#0436# => romdata <= X"13C09F46";
    when 16#0437# => romdata <= X"8DC97FC0";
    when 16#0438# => romdata <= X"E5DD057A";
    when 16#0439# => romdata <= X"8A035576";
    when 16#043A# => romdata <= X"7B698F8A";
    when 16#043B# => romdata <= X"79BF0350";
    when 16#043C# => romdata <= X"C4200413";
    when 16#043D# => romdata <= X"A15E6591";
    when 16#043E# => romdata <= X"DE70A1B5";
    when 16#043F# => romdata <= X"02E19FF5";
    when 16#0440# => romdata <= X"15C3DF36";
    when 16#0441# => romdata <= X"935974A4";
    when 16#0442# => romdata <= X"764895B9";
    when 16#0443# => romdata <= X"E3CA2626";
    when 16#0444# => romdata <= X"BD39B7AD";
    when 16#0445# => romdata <= X"B780AAF7";
    when 16#0446# => romdata <= X"E2E914E8";
    when 16#0447# => romdata <= X"04CA9230";
    when 16#0448# => romdata <= X"89A51F38";
    when 16#0449# => romdata <= X"76649C73";
    when 16#044A# => romdata <= X"CA3C2623";
    when 16#044B# => romdata <= X"A8C95D11";
    when 16#044C# => romdata <= X"EF4B3F94";
    when 16#044D# => romdata <= X"1E9772EB";
    when 16#044E# => romdata <= X"A1F47212";
    when 16#044F# => romdata <= X"C666F03F";
    when 16#0450# => romdata <= X"01509FF6";
    when 16#0451# => romdata <= X"99F74EDE";
    when 16#0452# => romdata <= X"27182B6E";
    when 16#0453# => romdata <= X"98AF49D1";
    when 16#0454# => romdata <= X"BAACB41A";
    when 16#0455# => romdata <= X"328A8C34";
    when 16#0456# => romdata <= X"D6E8AA35";
    when 16#0457# => romdata <= X"53DA3962";
    when 16#0458# => romdata <= X"B27B0414";
    when 16#0459# => romdata <= X"95F26932";
    when 16#045A# => romdata <= X"8B6BFB4A";
    when 16#045B# => romdata <= X"385CBB11";
    when 16#045C# => romdata <= X"8953F3F0";
    when 16#045D# => romdata <= X"09920EC4";
    when 16#045E# => romdata <= X"C8590003";
    when 16#045F# => romdata <= X"290DD60A";
    when 16#0460# => romdata <= X"C89177BB";
    when 16#0461# => romdata <= X"8C4BF753";
    when 16#0462# => romdata <= X"CE723AEC";
    when 16#0463# => romdata <= X"A392B8D9";
    when 16#0464# => romdata <= X"E5E9E411";
    when 16#0465# => romdata <= X"3DD062F2";
    when 16#0466# => romdata <= X"94A77B6E";
    when 16#0467# => romdata <= X"A9A0477E";
    when 16#0468# => romdata <= X"697C04C7";
    when 16#0469# => romdata <= X"87CE78A9";
    when 16#046A# => romdata <= X"2C704409";
    when 16#046B# => romdata <= X"D37D37B6";
    when 16#046C# => romdata <= X"B3921286";
    when 16#046D# => romdata <= X"98D0D8D4";
    when 16#046E# => romdata <= X"CA101EB3";
    when 16#046F# => romdata <= X"8B92F467";
    when 16#0470# => romdata <= X"F0D86EFD";
    when 16#0471# => romdata <= X"8759A141";
    when 16#0472# => romdata <= X"62CAB55F";
    when 16#0473# => romdata <= X"8C457E82";
    when 16#0474# => romdata <= X"392790A5";
    when 16#0475# => romdata <= X"BDDC8DD2";
    when 16#0476# => romdata <= X"663944F8";
    when 16#0477# => romdata <= X"80C95EC0";
    when 16#0478# => romdata <= X"2FE5363B";
    when 16#0479# => romdata <= X"06462399";
    when 16#047A# => romdata <= X"4EE5D439";
    when 16#047B# => romdata <= X"6C0E44DE";
    when 16#047C# => romdata <= X"2A3D2258";
    when 16#047D# => romdata <= X"30BA6160";
    when 16#047E# => romdata <= X"270BCD11";
    when 16#047F# => romdata <= X"0A942B00";
    when 16#0480# => romdata <= X"92A0DEAB";
    when 16#0481# => romdata <= X"A9875D4A";
    when 16#0482# => romdata <= X"FAF99A24";
    when 16#0483# => romdata <= X"C1D5F10E";
    when 16#0484# => romdata <= X"BBE6DEF9";
    when 16#0485# => romdata <= X"CAE5B0C8";
    when 16#0486# => romdata <= X"5B2A0417";
    when 16#0487# => romdata <= X"C1CC5D1A";
    when 16#0488# => romdata <= X"5F71CD8F";
    when 16#0489# => romdata <= X"8A4B013C";
    when 16#048A# => romdata <= X"3F012C0A";
    when 16#048B# => romdata <= X"19EE4A23";
    when 16#048C# => romdata <= X"106CAB86";
    when 16#048D# => romdata <= X"62C5A2A9";
    when 16#048E# => romdata <= X"3A971D0B";
    when 16#048F# => romdata <= X"6E487FC0";
    when 16#0490# => romdata <= X"5BAF5C35";
    when 16#0491# => romdata <= X"5A9520C9";
    when 16#0492# => romdata <= X"148584CF";
    when 16#0493# => romdata <= X"ED3EDD0F";
    when 16#0494# => romdata <= X"38696E16";
    when 16#0495# => romdata <= X"1E64378C";
    when 16#0496# => romdata <= X"831C586D";
    when 16#0497# => romdata <= X"9178A0CE";
    when 16#0498# => romdata <= X"289A67F3";
    when 16#0499# => romdata <= X"3AE68C02";
    when 16#049A# => romdata <= X"A3CD138F";
    when 16#049B# => romdata <= X"A09DF1CA";
    when 16#049C# => romdata <= X"D01EFADF";
    when 16#049D# => romdata <= X"C8BF6F54";
    when 16#049E# => romdata <= X"07B79B18";
    when 16#049F# => romdata <= X"D09C8280";
    when 16#04A0# => romdata <= X"4736752D";
    when 16#04A1# => romdata <= X"08A1FE09";
    when 16#04A2# => romdata <= X"EB35F544";
    when 16#04A3# => romdata <= X"E9F797EA";
    when 16#04A4# => romdata <= X"36DB493B";
    when 16#04A5# => romdata <= X"A947AA82";
    when 16#04A6# => romdata <= X"513EB161";
    when 16#04A7# => romdata <= X"5A356B5A";
    when 16#04A8# => romdata <= X"A4308B0B";
    when 16#04A9# => romdata <= X"4183E070";
    when 16#04AA# => romdata <= X"EB494D62";
    when 16#04AB# => romdata <= X"8159D2D4";
    when 16#04AC# => romdata <= X"BC3CB110";
    when 16#04AD# => romdata <= X"AB0CCB2E";
    when 16#04AE# => romdata <= X"9E73B5B7";
    when 16#04AF# => romdata <= X"EB567187";
    when 16#04B0# => romdata <= X"621E72D9";
    when 16#04B1# => romdata <= X"9F1FB785";
    when 16#04B2# => romdata <= X"65917B28";
    when 16#04B3# => romdata <= X"464A5F29";
    when 16#04B4# => romdata <= X"DD8D6F98";
    when 16#04B5# => romdata <= X"B6ED7030";
    when 16#04B6# => romdata <= X"40A44B0A";
    when 16#04B7# => romdata <= X"CD97F150";
    when 16#04B8# => romdata <= X"49E009E8";
    when 16#04B9# => romdata <= X"533FDB0B";
    when 16#04BA# => romdata <= X"6DB2F258";
    when 16#04BB# => romdata <= X"2E6BBF81";
    when 16#04BC# => romdata <= X"D7B0EADC";
    when 16#04BD# => romdata <= X"8F402508";
    when 16#04BE# => romdata <= X"F6B8531A";
    when 16#04BF# => romdata <= X"D13FD1C5";
    when 16#04C0# => romdata <= X"5978A8A7";
    when 16#04C1# => romdata <= X"0DF4E053";
    when 16#04C2# => romdata <= X"DD475132";
    when 16#04C3# => romdata <= X"D348AE27";
    when 16#04C4# => romdata <= X"581370EC";
    when 16#04C5# => romdata <= X"14A3E0F9";
    when 16#04C6# => romdata <= X"6E0D70DA";
    when 16#04C7# => romdata <= X"4946DEEC";
    when 16#04C8# => romdata <= X"07600114";
    when 16#04C9# => romdata <= X"04FDC5B4";
    when 16#04CA# => romdata <= X"36CA7419";
    when 16#04CB# => romdata <= X"D05895F5";
    when 16#04CC# => romdata <= X"E0EAEEBC";
    when 16#04CD# => romdata <= X"88C74947";
    when 16#04CE# => romdata <= X"733BE991";
    when 16#04CF# => romdata <= X"9F18CE70";
    when 16#04D0# => romdata <= X"2887A6C4";
    when 16#04D1# => romdata <= X"DF7C1927";
    when 16#04D2# => romdata <= X"9B82FB64";
    when 16#04D3# => romdata <= X"6090822D";
    when 16#04D4# => romdata <= X"A9CD9C76";
    when 16#04D5# => romdata <= X"53F6B931";
    when 16#04D6# => romdata <= X"A337A28F";
    when 16#04D7# => romdata <= X"7A4A01DE";
    when 16#04D8# => romdata <= X"0CC0744F";
    when 16#04D9# => romdata <= X"22961045";
    when 16#04DA# => romdata <= X"F8EF8D4B";
    when 16#04DB# => romdata <= X"30B07E5E";
    when 16#04DC# => romdata <= X"DF5FA944";
    when 16#04DD# => romdata <= X"EDCFB984";
    when 16#04DE# => romdata <= X"1A9088AE";
    when 16#04DF# => romdata <= X"82444FCB";
    when 16#04E0# => romdata <= X"6E90B0E9";
    when 16#04E1# => romdata <= X"C567A80E";
    when 16#04E2# => romdata <= X"8C42EC71";
    when 16#04E3# => romdata <= X"3D78132F";
    when 16#04E4# => romdata <= X"37AD1D25";
    when 16#04E5# => romdata <= X"92C31C93";
    when 16#04E6# => romdata <= X"D2EAEFF3";
    when 16#04E7# => romdata <= X"8AD94E5C";
    when 16#04E8# => romdata <= X"0D94F949";
    when 16#04E9# => romdata <= X"F47B88B0";
    when 16#04EA# => romdata <= X"3BC1EA4E";
    when 16#04EB# => romdata <= X"5EC9C7D9";
    when 16#04EC# => romdata <= X"DF19ED20";
    when 16#04ED# => romdata <= X"8B8E44FF";
    when 16#04EE# => romdata <= X"DEB0B625";
    when 16#04EF# => romdata <= X"F633C7DB";
    when 16#04F0# => romdata <= X"1C826AA9";
    when 16#04F1# => romdata <= X"E1C1309E";
    when 16#04F2# => romdata <= X"5B14A0DD";
    when 16#04F3# => romdata <= X"DB79714D";
    when 16#04F4# => romdata <= X"FDCB5222";
    when 16#04F5# => romdata <= X"1CEAD7E8";
    when 16#04F6# => romdata <= X"A140DF78";
    when 16#04F7# => romdata <= X"06F12715";
    when 16#04F8# => romdata <= X"6478AFBE";
    when 16#04F9# => romdata <= X"E922B8EC";
    when 16#04FA# => romdata <= X"F322D66B";
    when 16#04FB# => romdata <= X"48BEC434";
    when 16#04FC# => romdata <= X"299BBB36";
    when 16#04FD# => romdata <= X"B3BD9030";
    when 16#04FE# => romdata <= X"467B7F2E";
    when 16#04FF# => romdata <= X"BBDF3580";
    when 16#0500# => romdata <= X"AFA7FBAC";
    when 16#0501# => romdata <= X"93326D0C";
    when 16#0502# => romdata <= X"36A38883";
    when 16#0503# => romdata <= X"1B99DF4D";
    when 16#0504# => romdata <= X"527BCE7C";
    when 16#0505# => romdata <= X"9070F7B4";
    when 16#0506# => romdata <= X"6B5FFCDE";
    when 16#0507# => romdata <= X"B0738480";
    when 16#0508# => romdata <= X"1AE5F86A";
    when 16#0509# => romdata <= X"89934DE2";
    when 16#050A# => romdata <= X"3DFE2C1A";
    when 16#050B# => romdata <= X"D117797D";
    when 16#050C# => romdata <= X"4FA1BBA6";
    when 16#050D# => romdata <= X"175823B4";
    when 16#050E# => romdata <= X"1166DBE9";
    when 16#050F# => romdata <= X"D126F17B";
    when 16#0510# => romdata <= X"3761E2C3";
    when 16#0511# => romdata <= X"52AB396A";
    when 16#0512# => romdata <= X"5A9CCEA4";
    when 16#0513# => romdata <= X"2A5E9EA1";
    when 16#0514# => romdata <= X"BE3497C0";
    when 16#0515# => romdata <= X"A5BA9121";
    when 16#0516# => romdata <= X"DB97F641";
    when 16#0517# => romdata <= X"59AAC78E";
    when 16#0518# => romdata <= X"62D7DEFF";
    when 16#0519# => romdata <= X"3BF4CF73";
    when 16#051A# => romdata <= X"F8CFBE04";
    when 16#051B# => romdata <= X"5C9D39E4";
    when 16#051C# => romdata <= X"1D5D208D";
    when 16#051D# => romdata <= X"CC4B47CA";
    when 16#051E# => romdata <= X"27E900C3";
    when 16#051F# => romdata <= X"CD8FD140";
    when 16#0520# => romdata <= X"8DC5E0F5";
    when 16#0521# => romdata <= X"114F2FE6";
    when 16#0522# => romdata <= X"5817D37C";
    when 16#0523# => romdata <= X"D1452C49";
    when 16#0524# => romdata <= X"67ACAA21";
    when 16#0525# => romdata <= X"19FB8D60";
    when 16#0526# => romdata <= X"E5E2FD8A";
    when 16#0527# => romdata <= X"820D0AAD";
    when 16#0528# => romdata <= X"D88B94D4";
    when 16#0529# => romdata <= X"0435C095";
    when 16#052A# => romdata <= X"568AE639";
    when 16#052B# => romdata <= X"4D3B97C8";
    when 16#052C# => romdata <= X"35BA868A";
    when 16#052D# => romdata <= X"83083316";
    when 16#052E# => romdata <= X"C49C75D3";
    when 16#052F# => romdata <= X"6EFDD851";
    when 16#0530# => romdata <= X"65BE74A4";
    when 16#0531# => romdata <= X"F2B2D212";
    when 16#0532# => romdata <= X"95EBCE08";
    when 16#0533# => romdata <= X"5D9C4A47";
    when 16#0534# => romdata <= X"58FDD9CF";
    when 16#0535# => romdata <= X"71B97FDF";
    when 16#0536# => romdata <= X"34B7B63A";
    when 16#0537# => romdata <= X"5E9691DB";
    when 16#0538# => romdata <= X"DAB834D8";
    when 16#0539# => romdata <= X"7D5B52CA";
    when 16#053A# => romdata <= X"9A53032F";
    when 16#053B# => romdata <= X"FE821398";
    when 16#053C# => romdata <= X"616EA926";
    when 16#053D# => romdata <= X"25C2DB63";
    when 16#053E# => romdata <= X"3E379119";
    when 16#053F# => romdata <= X"87083A3B";
    when 16#0540# => romdata <= X"49A86FC5";
    when 16#0541# => romdata <= X"62FB1264";
    when 16#0542# => romdata <= X"A75643A5";
    when 16#0543# => romdata <= X"FB6E9716";
    when 16#0544# => romdata <= X"2E16ACCE";
    when 16#0545# => romdata <= X"353227FE";
    when 16#0546# => romdata <= X"61A859E0";
    when 16#0547# => romdata <= X"94C2359B";
    when 16#0548# => romdata <= X"C4645946";
    when 16#0549# => romdata <= X"AD12AE5C";
    when 16#054A# => romdata <= X"39C70F59";
    when 16#054B# => romdata <= X"EA7B597A";
    when 16#054C# => romdata <= X"9B3372C2";
    when 16#054D# => romdata <= X"3AA57814";
    when 16#054E# => romdata <= X"6781A611";
    when 16#054F# => romdata <= X"63C92816";
    when 16#0550# => romdata <= X"627DD9C4";
    when 16#0551# => romdata <= X"BF178808";
    when 16#0552# => romdata <= X"7821F9F5";
    when 16#0553# => romdata <= X"D41B75A0";
    when 16#0554# => romdata <= X"F251B06B";
    when 16#0555# => romdata <= X"BD3E29AB";
    when 16#0556# => romdata <= X"D41E72A1";
    when 16#0557# => romdata <= X"D48323D2";
    when 16#0558# => romdata <= X"4E2AD6F1";
    when 16#0559# => romdata <= X"1C2D4967";
    when 16#055A# => romdata <= X"8CC04FCF";
    when 16#055B# => romdata <= X"6B0EFD33";
    when 16#055C# => romdata <= X"BE6DDCD4";
    when 16#055D# => romdata <= X"44F5CA02";
    when 16#055E# => romdata <= X"FE158112";
    when 16#055F# => romdata <= X"631F782C";
    when 16#0560# => romdata <= X"A7B0C5F3";
    when 16#0561# => romdata <= X"607ED807";
    when 16#0562# => romdata <= X"495BF8E8";
    when 16#0563# => romdata <= X"2C5EA51A";
    when 16#0564# => romdata <= X"922FE28C";
    when 16#0565# => romdata <= X"8168D984";
    when 16#0566# => romdata <= X"4859E7A3";
    when 16#0567# => romdata <= X"EE3038C5";
    when 16#0568# => romdata <= X"D1D4BB4B";
    when 16#0569# => romdata <= X"13406C34";
    when 16#056A# => romdata <= X"0894DF46";
    when 16#056B# => romdata <= X"40683673";
    when 16#056C# => romdata <= X"9E31D010";
    when 16#056D# => romdata <= X"82BC8448";
    when 16#056E# => romdata <= X"9592DA0E";
    when 16#056F# => romdata <= X"985630CE";
    when 16#0570# => romdata <= X"C40702A3";
    when 16#0571# => romdata <= X"6DDC301B";
    when 16#0572# => romdata <= X"3AE1E810";
    when 16#0573# => romdata <= X"1786FEDB";
    when 16#0574# => romdata <= X"F752F9E1";
    when 16#0575# => romdata <= X"75287C23";
    when 16#0576# => romdata <= X"9C18FC25";
    when 16#0577# => romdata <= X"795BCB47";
    when 16#0578# => romdata <= X"9DEF59C5";
    when 16#0579# => romdata <= X"8C373313";
    when 16#057A# => romdata <= X"C02A1BC5";
    when 16#057B# => romdata <= X"F16355E2";
    when 16#057C# => romdata <= X"B50EFB58";
    when 16#057D# => romdata <= X"85567086";
    when 16#057E# => romdata <= X"8728B902";
    when 16#057F# => romdata <= X"653ED800";
    when 16#0580# => romdata <= X"943CAEB6";
    when 16#0581# => romdata <= X"80AA3E63";
    when 16#0582# => romdata <= X"0755DF32";
    when 16#0583# => romdata <= X"F406F403";
    when 16#0584# => romdata <= X"D7AF5E48";
    when 16#0585# => romdata <= X"A710274D";
    when 16#0586# => romdata <= X"3887A7AA";
    when 16#0587# => romdata <= X"C8EA6744";
    when 16#0588# => romdata <= X"B889F2E0";
    when 16#0589# => romdata <= X"CD2033DE";
    when 16#058A# => romdata <= X"C0B434A9";
    when 16#058B# => romdata <= X"591254A0";
    when 16#058C# => romdata <= X"AA68C5C9";
    when 16#058D# => romdata <= X"BF11D357";
    when 16#058E# => romdata <= X"65E86B43";
    when 16#058F# => romdata <= X"7497D84E";
    when 16#0590# => romdata <= X"5DCBBC0C";
    when 16#0591# => romdata <= X"0C580CE9";
    when 16#0592# => romdata <= X"BC50EC63";
    when 16#0593# => romdata <= X"82AD74DB";
    when 16#0594# => romdata <= X"02C2C233";
    when 16#0595# => romdata <= X"B7BB0751";
    when 16#0596# => romdata <= X"7D480562";
    when 16#0597# => romdata <= X"26C505AB";
    when 16#0598# => romdata <= X"F2DD244F";
    when 16#0599# => romdata <= X"6BBAA233";
    when 16#059A# => romdata <= X"13D57055";
    when 16#059B# => romdata <= X"8B065E42";
    when 16#059C# => romdata <= X"32776807";
    when 16#059D# => romdata <= X"8EFDB53D";
    when 16#059E# => romdata <= X"C465DA03";
    when 16#059F# => romdata <= X"8E3B216D";
    when 16#05A0# => romdata <= X"990EE951";
    when 16#05A1# => romdata <= X"B3E13D3C";
    when 16#05A2# => romdata <= X"1CD55999";
    when 16#05A3# => romdata <= X"8F77BCDC";
    when 16#05A4# => romdata <= X"D2B9522B";
    when 16#05A5# => romdata <= X"6F1DC5E1";
    when 16#05A6# => romdata <= X"2C912EAE";
    when 16#05A7# => romdata <= X"F574AFD6";
    when 16#05A8# => romdata <= X"9C251F9B";
    when 16#05A9# => romdata <= X"2532501A";
    when 16#05AA# => romdata <= X"B9F4B3B2";
    when 16#05AB# => romdata <= X"223D0F89";
    when 16#05AC# => romdata <= X"20BD562B";
    when 16#05AD# => romdata <= X"0D358A14";
    when 16#05AE# => romdata <= X"AB0D196D";
    when 16#05AF# => romdata <= X"F6337D1C";
    when 16#05B0# => romdata <= X"96CDB47A";
    when 16#05B1# => romdata <= X"FEC6F81D";
    when 16#05B2# => romdata <= X"ED4B5773";
    when 16#05B3# => romdata <= X"864DA32F";
    when 16#05B4# => romdata <= X"CCD06B9A";
    when 16#05B5# => romdata <= X"C53C122B";
    when 16#05B6# => romdata <= X"2C6327E6";
    when 16#05B7# => romdata <= X"E5EFE227";
    when 16#05B8# => romdata <= X"DE4893FF";
    when 16#05B9# => romdata <= X"15BBB225";
    when 16#05BA# => romdata <= X"7FAEA836";
    when 16#05BB# => romdata <= X"E99676EE";
    when 16#05BC# => romdata <= X"32BF6FC1";
    when 16#05BD# => romdata <= X"4D4F56EA";
    when 16#05BE# => romdata <= X"191B8A38";
    when 16#05BF# => romdata <= X"70374A08";
    when 16#05C0# => romdata <= X"67C49EB0";
    when 16#05C1# => romdata <= X"015D1C6D";
    when 16#05C2# => romdata <= X"07B87A36";
    when 16#05C3# => romdata <= X"BFDD1DCE";
    when 16#05C4# => romdata <= X"F20EA7B8";
    when 16#05C5# => romdata <= X"0D997CBE";
    when 16#05C6# => romdata <= X"2D83EB56";
    when 16#05C7# => romdata <= X"30F2EE6F";
    when 16#05C8# => romdata <= X"73B0D507";
    when 16#05C9# => romdata <= X"00C89E4F";
    when 16#05CA# => romdata <= X"32438F55";
    when 16#05CB# => romdata <= X"41360683";
    when 16#05CC# => romdata <= X"DF11DA6E";
    when 16#05CD# => romdata <= X"7A3C1E7D";
    when 16#05CE# => romdata <= X"B2A87800";
    when 16#05CF# => romdata <= X"D9245BF0";
    when 16#05D0# => romdata <= X"4278C990";
    when 16#05D1# => romdata <= X"A8DC9CD8";
    when 16#05D2# => romdata <= X"6DEF39CB";
    when 16#05D3# => romdata <= X"C6D4BC00";
    when 16#05D4# => romdata <= X"FF13BBE1";
    when 16#05D5# => romdata <= X"32F9D866";
    when 16#05D6# => romdata <= X"81A8913B";
    when 16#05D7# => romdata <= X"E787CFC6";
    when 16#05D8# => romdata <= X"9C353048";
    when 16#05D9# => romdata <= X"24788716";
    when 16#05DA# => romdata <= X"D52DC74C";
    when 16#05DB# => romdata <= X"EA399E06";
    when 16#05DC# => romdata <= X"DE624178";
    when 16#05DD# => romdata <= X"0447C74D";
    when 16#05DE# => romdata <= X"A8E94713";
    when 16#05DF# => romdata <= X"4D8B2FAA";
    when 16#05E0# => romdata <= X"9648D6D5";
    when 16#05E1# => romdata <= X"F34C9D60";
    when 16#05E2# => romdata <= X"AE5973B5";
    when 16#05E3# => romdata <= X"BB018779";
    when 16#05E4# => romdata <= X"6D589C8F";
    when 16#05E5# => romdata <= X"DDD76756";
    when 16#05E6# => romdata <= X"71F28C04";
    when 16#05E7# => romdata <= X"AC1038D0";
    when 16#05E8# => romdata <= X"92519806";
    when 16#05E9# => romdata <= X"83CB712F";
    when 16#05EA# => romdata <= X"694D7C5B";
    when 16#05EB# => romdata <= X"0D5B1DE8";
    when 16#05EC# => romdata <= X"6CD10EAC";
    when 16#05ED# => romdata <= X"4EA04A55";
    when 16#05EE# => romdata <= X"BA8803D7";
    when 16#05EF# => romdata <= X"8249BEF5";
    when 16#05F0# => romdata <= X"16D38067";
    when 16#05F1# => romdata <= X"890105A2";
    when 16#05F2# => romdata <= X"3212E728";
    when 16#05F3# => romdata <= X"79FA267A";
    when 16#05F4# => romdata <= X"8B4F0455";
    when 16#05F5# => romdata <= X"A81F17CF";
    when 16#05F6# => romdata <= X"D3E5DDC5";
    when 16#05F7# => romdata <= X"5E5D4FE0";
    when 16#05F8# => romdata <= X"0F83E186";
    when 16#05F9# => romdata <= X"26C676DA";
    when 16#05FA# => romdata <= X"F00E6AAF";
    when 16#05FB# => romdata <= X"CC23D209";
    when 16#05FC# => romdata <= X"DEE0B0FC";
    when 16#05FD# => romdata <= X"6C2AE4DE";
    when 16#05FE# => romdata <= X"161D1301";
    when 16#05FF# => romdata <= X"7ADB5D80";
    when 16#0600# => romdata <= X"E5E70E78";
    when 16#0601# => romdata <= X"37D09441";
    when 16#0602# => romdata <= X"6558C044";
    when 16#0603# => romdata <= X"D758383E";
    when 16#0604# => romdata <= X"DF5755C8";
    when 16#0605# => romdata <= X"0921218A";
    when 16#0606# => romdata <= X"BE76E51F";
    when 16#0607# => romdata <= X"B93249E2";
    when 16#0608# => romdata <= X"11A38FE6";
    when 16#0609# => romdata <= X"D07A7DFD";
    when 16#060A# => romdata <= X"2263E6E3";
    when 16#060B# => romdata <= X"D8DA0F92";
    when 16#060C# => romdata <= X"1A06A606";
    when 16#060D# => romdata <= X"B804DE7A";
    when 16#060E# => romdata <= X"C3FD097E";
    when 16#060F# => romdata <= X"5F96EFCC";
    when 16#0610# => romdata <= X"0F544D62";
    when 16#0611# => romdata <= X"3FD6F43F";
    when 16#0612# => romdata <= X"B88CEA7C";
    when 16#0613# => romdata <= X"341E901C";
    when 16#0614# => romdata <= X"D47A7E24";
    when 16#0615# => romdata <= X"AB141E99";
    when 16#0616# => romdata <= X"8FE41CA8";
    when 16#0617# => romdata <= X"7CD6CE8C";
    when 16#0618# => romdata <= X"1870D9AB";
    when 16#0619# => romdata <= X"B6503BF7";
    when 16#061A# => romdata <= X"E8B65908";
    when 16#061B# => romdata <= X"4BAF2237";
    when 16#061C# => romdata <= X"DFC94F35";
    when 16#061D# => romdata <= X"C9884C7F";
    when 16#061E# => romdata <= X"44B87120";
    when 16#061F# => romdata <= X"BFCB2986";
    when 16#0620# => romdata <= X"96E613C1";
    when 16#0621# => romdata <= X"656AC489";
    when 16#0622# => romdata <= X"9781A948";
    when 16#0623# => romdata <= X"69EC603B";
    when 16#0624# => romdata <= X"4D386653";
    when 16#0625# => romdata <= X"37CA8593";
    when 16#0626# => romdata <= X"AAC83AD8";
    when 16#0627# => romdata <= X"BECE1030";
    when 16#0628# => romdata <= X"2E4B4694";
    when 16#0629# => romdata <= X"237E96CC";
    when 16#062A# => romdata <= X"D3AD9CD5";
    when 16#062B# => romdata <= X"F8EC039A";
    when 16#062C# => romdata <= X"1D1A4210";
    when 16#062D# => romdata <= X"71637140";
    when 16#062E# => romdata <= X"4C5C3FF3";
    when 16#062F# => romdata <= X"75CB3A33";
    when 16#0630# => romdata <= X"559B1C1A";
    when 16#0631# => romdata <= X"239F2E44";
    when 16#0632# => romdata <= X"2C8EB033";
    when 16#0633# => romdata <= X"501BB290";
    when 16#0634# => romdata <= X"434BE734";
    when 16#0635# => romdata <= X"89F71696";
    when 16#0636# => romdata <= X"53939894";
    when 16#0637# => romdata <= X"22CF4D57";
    when 16#0638# => romdata <= X"E5B4F3C7";
    when 16#0639# => romdata <= X"6AF3C5E8";
    when 16#063A# => romdata <= X"999E6180";
    when 16#063B# => romdata <= X"5134B9D7";
    when 16#063C# => romdata <= X"C40BFB59";
    when 16#063D# => romdata <= X"D0D0FD30";
    when 16#063E# => romdata <= X"F98567E6";
    when 16#063F# => romdata <= X"6D6148D6";
    when 16#0640# => romdata <= X"AA64F74A";
    when 16#0641# => romdata <= X"22C50AE4";
    when 16#0642# => romdata <= X"9D6B1ECC";
    when 16#0643# => romdata <= X"6BB5A002";
    when 16#0644# => romdata <= X"ABF38FF2";
    when 16#0645# => romdata <= X"E2436766";
    when 16#0646# => romdata <= X"B86BDDE7";
    when 16#0647# => romdata <= X"D95DD6E0";
    when 16#0648# => romdata <= X"2AB0FF06";
    when 16#0649# => romdata <= X"E7BC22CE";
    when 16#064A# => romdata <= X"C98D55AA";
    when 16#064B# => romdata <= X"2BC4D7B9";
    when 16#064C# => romdata <= X"1C36B2FF";
    when 16#064D# => romdata <= X"9F525A74";
    when 16#064E# => romdata <= X"423498D5";
    when 16#064F# => romdata <= X"48318509";
    when 16#0650# => romdata <= X"320FCCBC";
    when 16#0651# => romdata <= X"A582A6C2";
    when 16#0652# => romdata <= X"996AF653";
    when 16#0653# => romdata <= X"8422FF0D";
    when 16#0654# => romdata <= X"F060C0BC";
    when 16#0655# => romdata <= X"7356B085";
    when 16#0656# => romdata <= X"0A139AC3";
    when 16#0657# => romdata <= X"91433812";
    when 16#0658# => romdata <= X"7B786F4B";
    when 16#0659# => romdata <= X"C58CEB60";
    when 16#065A# => romdata <= X"64DA8813";
    when 16#065B# => romdata <= X"76A147DF";
    when 16#065C# => romdata <= X"F53C6700";
    when 16#065D# => romdata <= X"BD13316A";
    when 16#065E# => romdata <= X"5874A75D";
    when 16#065F# => romdata <= X"7B9713DF";
    when 16#0660# => romdata <= X"54FBB393";
    when 16#0661# => romdata <= X"BAFAAD7F";
    when 16#0662# => romdata <= X"7B0710C0";
    when 16#0663# => romdata <= X"49A0B6A8";
    when 16#0664# => romdata <= X"B76A9956";
    when 16#0665# => romdata <= X"BF6185BA";
    when 16#0666# => romdata <= X"39D9C347";
    when 16#0667# => romdata <= X"D179FBB9";
    when 16#0668# => romdata <= X"7D4FED68";
    when 16#0669# => romdata <= X"F47DB5AC";
    when 16#066A# => romdata <= X"8E0D4012";
    when 16#066B# => romdata <= X"2EA51C4A";
    when 16#066C# => romdata <= X"1F88D231";
    when 16#066D# => romdata <= X"53DF651A";
    when 16#066E# => romdata <= X"180C2AD4";
    when 16#066F# => romdata <= X"56ABD7F8";
    when 16#0670# => romdata <= X"51B65B22";
    when 16#0671# => romdata <= X"0A72BA48";
    when 16#0672# => romdata <= X"FAD04363";
    when 16#0673# => romdata <= X"32E4EE7E";
    when 16#0674# => romdata <= X"DC554B7D";
    when 16#0675# => romdata <= X"75481EE0";
    when 16#0676# => romdata <= X"5C3D3453";
    when 16#0677# => romdata <= X"D760E909";
    when 16#0678# => romdata <= X"9DD27B32";
    when 16#0679# => romdata <= X"4DD84C0C";
    when 16#067A# => romdata <= X"0C4DEC4C";
    when 16#067B# => romdata <= X"674D2528";
    when 16#067C# => romdata <= X"4B16410F";
    when 16#067D# => romdata <= X"959FBD09";
    when 16#067E# => romdata <= X"D9DF09CE";
    when 16#067F# => romdata <= X"875601E0";
    when 16#0680# => romdata <= X"BFDBC82A";
    when 16#0681# => romdata <= X"CB4FBCD5";
    when 16#0682# => romdata <= X"A90C5967";
    when 16#0683# => romdata <= X"EB2FED59";
    when 16#0684# => romdata <= X"7A02607F";
    when 16#0685# => romdata <= X"42600212";
    when 16#0686# => romdata <= X"8AF4B389";
    when 16#0687# => romdata <= X"42C85AF4";
    when 16#0688# => romdata <= X"472B3CBF";
    when 16#0689# => romdata <= X"3B183F24";
    when 16#068A# => romdata <= X"0E049B25";
    when 16#068B# => romdata <= X"1713740A";
    when 16#068C# => romdata <= X"31117F10";
    when 16#068D# => romdata <= X"8936631F";
    when 16#068E# => romdata <= X"D0F11C5F";
    when 16#068F# => romdata <= X"79325BD6";
    when 16#0690# => romdata <= X"677A2C2B";
    when 16#0691# => romdata <= X"242965AE";
    when 16#0692# => romdata <= X"FC147D93";
    when 16#0693# => romdata <= X"358730AA";
    when 16#0694# => romdata <= X"78249120";
    when 16#0695# => romdata <= X"9CBE6009";
    when 16#0696# => romdata <= X"76F56030";
    when 16#0697# => romdata <= X"753CC979";
    when 16#0698# => romdata <= X"C240A196";
    when 16#0699# => romdata <= X"647CD9EA";
    when 16#069A# => romdata <= X"B1DD0380";
    when 16#069B# => romdata <= X"E59BC790";
    when 16#069C# => romdata <= X"5EF740C3";
    when 16#069D# => romdata <= X"411AD9DD";
    when 16#069E# => romdata <= X"72027D0D";
    when 16#069F# => romdata <= X"3DD6DEB0";
    when 16#06A0# => romdata <= X"F5F3C18F";
    when 16#06A1# => romdata <= X"6D6F7BC5";
    when 16#06A2# => romdata <= X"9B758E7E";
    when 16#06A3# => romdata <= X"262937B4";
    when 16#06A4# => romdata <= X"599B3856";
    when 16#06A5# => romdata <= X"7C147ED2";
    when 16#06A6# => romdata <= X"689BA2CF";
    when 16#06A7# => romdata <= X"23736CAF";
    when 16#06A8# => romdata <= X"55B69258";
    when 16#06A9# => romdata <= X"27E2B70E";
    when 16#06AA# => romdata <= X"47D3813C";
    when 16#06AB# => romdata <= X"94C85298";
    when 16#06AC# => romdata <= X"BD6B49C9";
    when 16#06AD# => romdata <= X"7B5D0221";
    when 16#06AE# => romdata <= X"BE9E3164";
    when 16#06AF# => romdata <= X"B6FA3D95";
    when 16#06B0# => romdata <= X"AECF53AF";
    when 16#06B1# => romdata <= X"17096609";
    when 16#06B2# => romdata <= X"0F19A69E";
    when 16#06B3# => romdata <= X"75F188BD";
    when 16#06B4# => romdata <= X"2556B4E8";
    when 16#06B5# => romdata <= X"FA7DC4AC";
    when 16#06B6# => romdata <= X"6C34F542";
    when 16#06B7# => romdata <= X"97C06C2A";
    when 16#06B8# => romdata <= X"96DD1C45";
    when 16#06B9# => romdata <= X"B42E6175";
    when 16#06BA# => romdata <= X"B5E87845";
    when 16#06BB# => romdata <= X"68F7FEF0";
    when 16#06BC# => romdata <= X"B6C124C5";
    when 16#06BD# => romdata <= X"019CB577";
    when 16#06BE# => romdata <= X"B374941E";
    when 16#06BF# => romdata <= X"8515CCFC";
    when 16#06C0# => romdata <= X"21F46D18";
    when 16#06C1# => romdata <= X"8BDD2C22";
    when 16#06C2# => romdata <= X"84C68887";
    when 16#06C3# => romdata <= X"9A5BEC50";
    when 16#06C4# => romdata <= X"CCB97FAE";
    when 16#06C5# => romdata <= X"E1F75580";
    when 16#06C6# => romdata <= X"577498D5";
    when 16#06C7# => romdata <= X"09D3DE16";
    when 16#06C8# => romdata <= X"1BE216C8";
    when 16#06C9# => romdata <= X"73B29E17";
    when 16#06CA# => romdata <= X"8CE17DCA";
    when 16#06CB# => romdata <= X"CC5E9E22";
    when 16#06CC# => romdata <= X"24D05ECC";
    when 16#06CD# => romdata <= X"842FBEAB";
    when 16#06CE# => romdata <= X"82A75AAA";
    when 16#06CF# => romdata <= X"20769FD8";
    when 16#06D0# => romdata <= X"1131CFB6";
    when 16#06D1# => romdata <= X"9D5E3540";
    when 16#06D2# => romdata <= X"9273CA10";
    when 16#06D3# => romdata <= X"6FFB27F6";
    when 16#06D4# => romdata <= X"3FF997CB";
    when 16#06D5# => romdata <= X"500F161F";
    when 16#06D6# => romdata <= X"6DD3A8BF";
    when 16#06D7# => romdata <= X"A5719F00";
    when 16#06D8# => romdata <= X"4EC17860";
    when 16#06D9# => romdata <= X"152D3290";
    when 16#06DA# => romdata <= X"951678A1";
    when 16#06DB# => romdata <= X"31E4F3D3";
    when 16#06DC# => romdata <= X"AB34CFFC";
    when 16#06DD# => romdata <= X"AB2967ED";
    when 16#06DE# => romdata <= X"9D8F1BB9";
    when 16#06DF# => romdata <= X"87950306";
    when 16#06E0# => romdata <= X"BD28751D";
    when 16#06E1# => romdata <= X"2AEAB05F";
    when 16#06E2# => romdata <= X"071B0857";
    when 16#06E3# => romdata <= X"4EFCA01E";
    when 16#06E4# => romdata <= X"5386E04F";
    when 16#06E5# => romdata <= X"727BF413";
    when 16#06E6# => romdata <= X"A8279E93";
    when 16#06E7# => romdata <= X"92EFB64D";
    when 16#06E8# => romdata <= X"9AEE0087";
    when 16#06E9# => romdata <= X"7C76C81E";
    when 16#06EA# => romdata <= X"BC861E2B";
    when 16#06EB# => romdata <= X"484A2D35";
    when 16#06EC# => romdata <= X"E592A131";
    when 16#06ED# => romdata <= X"726CAE61";
    when 16#06EE# => romdata <= X"BC010B95";
    when 16#06EF# => romdata <= X"4721A82C";
    when 16#06F0# => romdata <= X"968CC6F3";
    when 16#06F1# => romdata <= X"84D9BBB9";
    when 16#06F2# => romdata <= X"9B4E8784";
    when 16#06F3# => romdata <= X"6D10B94E";
    when 16#06F4# => romdata <= X"E31F6484";
    when 16#06F5# => romdata <= X"6A5834DF";
    when 16#06F6# => romdata <= X"73A67A26";
    when 16#06F7# => romdata <= X"7B894B1C";
    when 16#06F8# => romdata <= X"06242D75";
    when 16#06F9# => romdata <= X"0F15F3E1";
    when 16#06FA# => romdata <= X"E850A11C";
    when 16#06FB# => romdata <= X"B2E2B161";
    when 16#06FC# => romdata <= X"55008F91";
    when 16#06FD# => romdata <= X"493AB3BC";
    when 16#06FE# => romdata <= X"77CF9BE5";
    when 16#06FF# => romdata <= X"6F9DB200";
    when 16#0700# => romdata <= X"D64F3D1C";
    when 16#0701# => romdata <= X"B54CDB91";
    when 16#0702# => romdata <= X"43D9E701";
    when 16#0703# => romdata <= X"BD313779";
    when 16#0704# => romdata <= X"C09DA064";
    when 16#0705# => romdata <= X"D9A85674";
    when 16#0706# => romdata <= X"CCB53B0C";
    when 16#0707# => romdata <= X"5B4446C1";
    when 16#0708# => romdata <= X"22098961";
    when 16#0709# => romdata <= X"D5EFFD6A";
    when 16#070A# => romdata <= X"85537486";
    when 16#070B# => romdata <= X"D5EB26B5";
    when 16#070C# => romdata <= X"E18FFBFB";
    when 16#070D# => romdata <= X"8E6EF16C";
    when 16#070E# => romdata <= X"2DD2C02E";
    when 16#070F# => romdata <= X"C7C07DB1";
    when 16#0710# => romdata <= X"5CE33015";
    when 16#0711# => romdata <= X"A636E225";
    when 16#0712# => romdata <= X"F744C963";
    when 16#0713# => romdata <= X"BF0653A8";
    when 16#0714# => romdata <= X"9A48F1AF";
    when 16#0715# => romdata <= X"04819E27";
    when 16#0716# => romdata <= X"3A3AE1F5";
    when 16#0717# => romdata <= X"538AD574";
    when 16#0718# => romdata <= X"D553C5A0";
    when 16#0719# => romdata <= X"DEF47B55";
    when 16#071A# => romdata <= X"2957037B";
    when 16#071B# => romdata <= X"CA921970";
    when 16#071C# => romdata <= X"C76DDEF7";
    when 16#071D# => romdata <= X"4BA083ED";
    when 16#071E# => romdata <= X"55363760";
    when 16#071F# => romdata <= X"A6780612";
    when 16#0720# => romdata <= X"C075964B";
    when 16#0721# => romdata <= X"083B4F67";
    when 16#0722# => romdata <= X"4EA0012F";
    when 16#0723# => romdata <= X"D1DF09F0";
    when 16#0724# => romdata <= X"445CE75A";
    when 16#0725# => romdata <= X"69885209";
    when 16#0726# => romdata <= X"8206868A";
    when 16#0727# => romdata <= X"D8241E3B";
    when 16#0728# => romdata <= X"319FA8D2";
    when 16#0729# => romdata <= X"D86DE6E7";
    when 16#072A# => romdata <= X"631DF1AE";
    when 16#072B# => romdata <= X"B571F967";
    when 16#072C# => romdata <= X"6323E062";
    when 16#072D# => romdata <= X"7307F6D8";
    when 16#072E# => romdata <= X"F569536A";
    when 16#072F# => romdata <= X"758DE5ED";
    when 16#0730# => romdata <= X"AAEDF80F";
    when 16#0731# => romdata <= X"4335E3AF";
    when 16#0732# => romdata <= X"CAD07F70";
    when 16#0733# => romdata <= X"AAD5CD08";
    when 16#0734# => romdata <= X"CCA1E71B";
    when 16#0735# => romdata <= X"84D4D979";
    when 16#0736# => romdata <= X"31F924AC";
    when 16#0737# => romdata <= X"0010C081";
    when 16#0738# => romdata <= X"1972ACAA";
    when 16#0739# => romdata <= X"414B89FF";
    when 16#073A# => romdata <= X"F7917E65";
    when 16#073B# => romdata <= X"3BB31E9C";
    when 16#073C# => romdata <= X"DFC72595";
    when 16#073D# => romdata <= X"066C662C";
    when 16#073E# => romdata <= X"DB9BBC96";
    when 16#073F# => romdata <= X"152D46BF";
    when 16#0740# => romdata <= X"4E8C15A8";
    when 16#0741# => romdata <= X"D34809C4";
    when 16#0742# => romdata <= X"B9D79871";
    when 16#0743# => romdata <= X"BDF0B63F";
    when 16#0744# => romdata <= X"A294F2D6";
    when 16#0745# => romdata <= X"67624F6E";
    when 16#0746# => romdata <= X"0210CD40";
    when 16#0747# => romdata <= X"C92F1C03";
    when 16#0748# => romdata <= X"3C3D8BF0";
    when 16#0749# => romdata <= X"89EF85C4";
    when 16#074A# => romdata <= X"F571CA72";
    when 16#074B# => romdata <= X"7C71B231";
    when 16#074C# => romdata <= X"28A9B0FF";
    when 16#074D# => romdata <= X"D70CEA93";
    when 16#074E# => romdata <= X"C316FC4D";
    when 16#074F# => romdata <= X"69D79B08";
    when 16#0750# => romdata <= X"9107F292";
    when 16#0751# => romdata <= X"E03425B2";
    when 16#0752# => romdata <= X"552AF5AA";
    when 16#0753# => romdata <= X"18FDB9AF";
    when 16#0754# => romdata <= X"86EA1972";
    when 16#0755# => romdata <= X"B66B1276";
    when 16#0756# => romdata <= X"B0911943";
    when 16#0757# => romdata <= X"7E4DFB8F";
    when 16#0758# => romdata <= X"8E3972D9";
    when 16#0759# => romdata <= X"1A93816E";
    when 16#075A# => romdata <= X"BD7D8D71";
    when 16#075B# => romdata <= X"5CB47EFA";
    when 16#075C# => romdata <= X"742938B0";
    when 16#075D# => romdata <= X"B49FA27A";
    when 16#075E# => romdata <= X"291B0DEA";
    when 16#075F# => romdata <= X"1DF0B8F8";
    when 16#0760# => romdata <= X"78332103";
    when 16#0761# => romdata <= X"F45A9993";
    when 16#0762# => romdata <= X"6896181E";
    when 16#0763# => romdata <= X"51FF65C6";
    when 16#0764# => romdata <= X"995F57C2";
    when 16#0765# => romdata <= X"C54B8002";
    when 16#0766# => romdata <= X"DEFF54B0";
    when 16#0767# => romdata <= X"EB3131EE";
    when 16#0768# => romdata <= X"7D61030C";
    when 16#0769# => romdata <= X"33B5502C";
    when 16#076A# => romdata <= X"49CF398F";
    when 16#076B# => romdata <= X"EC4B7615";
    when 16#076C# => romdata <= X"D16FCEA3";
    when 16#076D# => romdata <= X"E8EA12BF";
    when 16#076E# => romdata <= X"B311D426";
    when 16#076F# => romdata <= X"331A0660";
    when 16#0770# => romdata <= X"6CA5A066";
    when 16#0771# => romdata <= X"707C4AF8";
    when 16#0772# => romdata <= X"D1048F1C";
    when 16#0773# => romdata <= X"A6065FBE";
    when 16#0774# => romdata <= X"506D06C6";
    when 16#0775# => romdata <= X"C00D5D25";
    when 16#0776# => romdata <= X"0E227265";
    when 16#0777# => romdata <= X"551867A6";
    when 16#0778# => romdata <= X"816F0515";
    when 16#0779# => romdata <= X"5FCBDE24";
    when 16#077A# => romdata <= X"D4AD115B";
    when 16#077B# => romdata <= X"DA98AFE0";
    when 16#077C# => romdata <= X"8B12A1F3";
    when 16#077D# => romdata <= X"2E7C2ADA";
    when 16#077E# => romdata <= X"801FFB78";
    when 16#077F# => romdata <= X"BA057260";
    when 16#0780# => romdata <= X"9D6AD988";
    when 16#0781# => romdata <= X"9EA02FC9";
    when 16#0782# => romdata <= X"A5894929";
    when 16#0783# => romdata <= X"0975DB0F";
    when 16#0784# => romdata <= X"512EB37C";
    when 16#0785# => romdata <= X"8156CC9F";
    when 16#0786# => romdata <= X"1242B9E4";
    when 16#0787# => romdata <= X"5F22CC1D";
    when 16#0788# => romdata <= X"6ED1CBCB";
    when 16#0789# => romdata <= X"6CB24581";
    when 16#078A# => romdata <= X"1CE72926";
    when 16#078B# => romdata <= X"1641FDF7";
    when 16#078C# => romdata <= X"A8F389BA";
    when 16#078D# => romdata <= X"FD7311B8";
    when 16#078E# => romdata <= X"BD689E02";
    when 16#078F# => romdata <= X"409F6E8C";
    when 16#0790# => romdata <= X"5202F466";
    when 16#0791# => romdata <= X"349EA466";
    when 16#0792# => romdata <= X"E5398B29";
    when 16#0793# => romdata <= X"C8CB126D";
    when 16#0794# => romdata <= X"9600D896";
    when 16#0795# => romdata <= X"97A07A69";
    when 16#0796# => romdata <= X"00FE8D95";
    when 16#0797# => romdata <= X"951903DA";
    when 16#0798# => romdata <= X"A3419839";
    when 16#0799# => romdata <= X"C2D9E35E";
    when 16#079A# => romdata <= X"9F4EABC0";
    when 16#079B# => romdata <= X"4C9006EA";
    when 16#079C# => romdata <= X"585F544C";
    when 16#079D# => romdata <= X"7163A33D";
    when 16#079E# => romdata <= X"7E78DE28";
    when 16#079F# => romdata <= X"256B7B89";
    when 16#07A0# => romdata <= X"78FE018C";
    when 16#07A1# => romdata <= X"B529F7F7";
    when 16#07A2# => romdata <= X"9BBF66DC";
    when 16#07A3# => romdata <= X"4F0DECE8";
    when 16#07A4# => romdata <= X"0AE3C2CD";
    when 16#07A5# => romdata <= X"479D78C4";
    when 16#07A6# => romdata <= X"480E4DE2";
    when 16#07A7# => romdata <= X"F06C70E5";
    when 16#07A8# => romdata <= X"FEBDFB4E";
    when 16#07A9# => romdata <= X"CAEDC2E7";
    when 16#07AA# => romdata <= X"BD891AD6";
    when 16#07AB# => romdata <= X"C91A7C24";
    when 16#07AC# => romdata <= X"46F1B13B";
    when 16#07AD# => romdata <= X"340B7160";
    when 16#07AE# => romdata <= X"782F6CC5";
    when 16#07AF# => romdata <= X"B45F9787";
    when 16#07B0# => romdata <= X"CF1B0985";
    when 16#07B1# => romdata <= X"202DDF02";
    when 16#07B2# => romdata <= X"EC552A6D";
    when 16#07B3# => romdata <= X"C41325FD";
    when 16#07B4# => romdata <= X"8D31A431";
    when 16#07B5# => romdata <= X"6C13C56F";
    when 16#07B6# => romdata <= X"7157134F";
    when 16#07B7# => romdata <= X"66E1D103";
    when 16#07B8# => romdata <= X"CC3AA7EB";
    when 16#07B9# => romdata <= X"951C9209";
    when 16#07BA# => romdata <= X"4EB4409E";
    when 16#07BB# => romdata <= X"6E7BC494";
    when 16#07BC# => romdata <= X"434FAD80";
    when 16#07BD# => romdata <= X"999D46D8";
    when 16#07BE# => romdata <= X"24A5A573";
    when 16#07BF# => romdata <= X"90599052";
    when 16#07C0# => romdata <= X"025F7DA4";
    when 16#07C1# => romdata <= X"838F7D16";
    when 16#07C2# => romdata <= X"A8DACDAF";
    when 16#07C3# => romdata <= X"A06D1755";
    when 16#07C4# => romdata <= X"46FADD1E";
    when 16#07C5# => romdata <= X"3F797526";
    when 16#07C6# => romdata <= X"5230F6C0";
    when 16#07C7# => romdata <= X"1B9C1FB1";
    when 16#07C8# => romdata <= X"B7AB1F2F";
    when 16#07C9# => romdata <= X"DD43A577";
    when 16#07CA# => romdata <= X"8E3C88FB";
    when 16#07CB# => romdata <= X"EA70575C";
    when 16#07CC# => romdata <= X"A26D94D2";
    when 16#07CD# => romdata <= X"49670E4D";
    when 16#07CE# => romdata <= X"9FF28EC6";
    when 16#07CF# => romdata <= X"7D158297";
    when 16#07D0# => romdata <= X"76D7BC67";
    when 16#07D1# => romdata <= X"54D2A2BB";
    when 16#07D2# => romdata <= X"01554E5F";
    when 16#07D3# => romdata <= X"F0C3FAD8";
    when 16#07D4# => romdata <= X"A1CB546E";
    when 16#07D5# => romdata <= X"8AD5E531";
    when 16#07D6# => romdata <= X"4103D086";
    when 16#07D7# => romdata <= X"D14ABD30";
    when 16#07D8# => romdata <= X"EA95DDC5";
    when 16#07D9# => romdata <= X"91C13D96";
    when 16#07DA# => romdata <= X"C1CC3F60";
    when 16#07DB# => romdata <= X"FD18D216";
    when 16#07DC# => romdata <= X"B67181B6";
    when 16#07DD# => romdata <= X"324AC09A";
    when 16#07DE# => romdata <= X"97C0C45E";
    when 16#07DF# => romdata <= X"50EE8380";
    when 16#07E0# => romdata <= X"ED42F6E0";
    when 16#07E1# => romdata <= X"43063937";
    when 16#07E2# => romdata <= X"3E7760C7";
    when 16#07E3# => romdata <= X"08248EE7";
    when 16#07E4# => romdata <= X"D74830E9";
    when 16#07E5# => romdata <= X"59411487";
    when 16#07E6# => romdata <= X"9748883F";
    when 16#07E7# => romdata <= X"247D056B";
    when 16#07E8# => romdata <= X"2BA94A0F";
    when 16#07E9# => romdata <= X"C54CECF6";
    when 16#07EA# => romdata <= X"F5C6AB4D";
    when 16#07EB# => romdata <= X"CB7CFC8C";
    when 16#07EC# => romdata <= X"224F40D8";
    when 16#07ED# => romdata <= X"86427504";
    when 16#07EE# => romdata <= X"233DDBED";
    when 16#07EF# => romdata <= X"CE160DEF";
    when 16#07F0# => romdata <= X"DFFD69EE";
    when 16#07F1# => romdata <= X"2B75746D";
    when 16#07F2# => romdata <= X"9CF71676";
    when 16#07F3# => romdata <= X"DC453FD0";
    when 16#07F4# => romdata <= X"1C315ACA";
    when 16#07F5# => romdata <= X"96373ED3";
    when 16#07F6# => romdata <= X"87B040BD";
    when 16#07F7# => romdata <= X"EBA7FF3C";
    when 16#07F8# => romdata <= X"E00D915F";
    when 16#07F9# => romdata <= X"90AE6E17";
    when 16#07FA# => romdata <= X"96971F80";
    when 16#07FB# => romdata <= X"52160154";
    when 16#07FC# => romdata <= X"E8986913";
    when 16#07FD# => romdata <= X"AD7BA291";
    when 16#07FE# => romdata <= X"188EC49A";
    when 16#07FF# => romdata <= X"60BE27C0";
    when 16#0800# => romdata <= X"B5184F7D";
    when 16#0801# => romdata <= X"580935AC";
    when 16#0802# => romdata <= X"FF18201C";
    when 16#0803# => romdata <= X"E8B5D54C";
    when 16#0804# => romdata <= X"D0A1CACF";
    when 16#0805# => romdata <= X"102FBC8A";
    when 16#0806# => romdata <= X"ADF391C4";
    when 16#0807# => romdata <= X"CA5807BA";
    when 16#0808# => romdata <= X"EEF4E5E4";
    when 16#0809# => romdata <= X"7F7459E7";
    when 16#080A# => romdata <= X"4485E48E";
    when 16#080B# => romdata <= X"0C42D27C";
    when 16#080C# => romdata <= X"ADE69707";
    when 16#080D# => romdata <= X"14FD97C0";
    when 16#080E# => romdata <= X"8F9592FD";
    when 16#080F# => romdata <= X"D387C859";
    when 16#0810# => romdata <= X"FC12C1CC";
    when 16#0811# => romdata <= X"CFC3EBF5";
    when 16#0812# => romdata <= X"10D66FBD";
    when 16#0813# => romdata <= X"8C448C25";
    when 16#0814# => romdata <= X"A322CC58";
    when 16#0815# => romdata <= X"87F94A55";
    when 16#0816# => romdata <= X"D48ECA36";
    when 16#0817# => romdata <= X"2C690F24";
    when 16#0818# => romdata <= X"833C3B03";
    when 16#0819# => romdata <= X"2A047D12";
    when 16#081A# => romdata <= X"BDA2ADC6";
    when 16#081B# => romdata <= X"824A1F6E";
    when 16#081C# => romdata <= X"A9320BED";
    when 16#081D# => romdata <= X"27968E9C";
    when 16#081E# => romdata <= X"FBDEC60D";
    when 16#081F# => romdata <= X"041EF538";
    when 16#0820# => romdata <= X"F1740C05";
    when 16#0821# => romdata <= X"19003FAA";
    when 16#0822# => romdata <= X"89CD4224";
    when 16#0823# => romdata <= X"293167E0";
    when 16#0824# => romdata <= X"5344998F";
    when 16#0825# => romdata <= X"D396EEF6";
    when 16#0826# => romdata <= X"18E8F547";
    when 16#0827# => romdata <= X"990BC06A";
    when 16#0828# => romdata <= X"8B76D0FD";
    when 16#0829# => romdata <= X"6FAC1328";
    when 16#082A# => romdata <= X"4601AB71";
    when 16#082B# => romdata <= X"91CEB813";
    when 16#082C# => romdata <= X"C46C45CE";
    when 16#082D# => romdata <= X"7B3FC09E";
    when 16#082E# => romdata <= X"DF08DAFE";
    when 16#082F# => romdata <= X"136BFBDD";
    when 16#0830# => romdata <= X"63E6CE7E";
    when 16#0831# => romdata <= X"4BCBB16C";
    when 16#0832# => romdata <= X"5DA68AC7";
    when 16#0833# => romdata <= X"1A1298FD";
    when 16#0834# => romdata <= X"27363349";
    when 16#0835# => romdata <= X"A261C2F2";
    when 16#0836# => romdata <= X"CA8CB799";
    when 16#0837# => romdata <= X"E8604ADF";
    when 16#0838# => romdata <= X"70092BDB";
    when 16#0839# => romdata <= X"D6A04CB8";
    when 16#083A# => romdata <= X"0568776A";
    when 16#083B# => romdata <= X"537AD171";
    when 16#083C# => romdata <= X"1891B251";
    when 16#083D# => romdata <= X"C74E42FC";
    when 16#083E# => romdata <= X"B095B23E";
    when 16#083F# => romdata <= X"EF70F167";
    when 16#0840# => romdata <= X"E8B4856B";
    when 16#0841# => romdata <= X"B7F92E3A";
    when 16#0842# => romdata <= X"43C79FF4";
    when 16#0843# => romdata <= X"437262DD";
    when 16#0844# => romdata <= X"70BAF9B1";
    when 16#0845# => romdata <= X"6CBF5F10";
    when 16#0846# => romdata <= X"D1AD7559";
    when 16#0847# => romdata <= X"AB0F8CEE";
    when 16#0848# => romdata <= X"1B9FAD05";
    when 16#0849# => romdata <= X"8E84FCC3";
    when 16#084A# => romdata <= X"42D9F0D9";
    when 16#084B# => romdata <= X"FBE4207D";
    when 16#084C# => romdata <= X"40E28141";
    when 16#084D# => romdata <= X"6506242C";
    when 16#084E# => romdata <= X"A1B8DAB2";
    when 16#084F# => romdata <= X"8DE88D2D";
    when 16#0850# => romdata <= X"00BA21AA";
    when 16#0851# => romdata <= X"7FDDC259";
    when 16#0852# => romdata <= X"40CB29F0";
    when 16#0853# => romdata <= X"2811F8DC";
    when 16#0854# => romdata <= X"6850A6A8";
    when 16#0855# => romdata <= X"7D72CA9F";
    when 16#0856# => romdata <= X"3476A736";
    when 16#0857# => romdata <= X"49FB4A25";
    when 16#0858# => romdata <= X"4B1204CC";
    when 16#0859# => romdata <= X"1261E7D5";
    when 16#085A# => romdata <= X"12BFE7B0";
    when 16#085B# => romdata <= X"D0091AD5";
    when 16#085C# => romdata <= X"CB0FBBB7";
    when 16#085D# => romdata <= X"65FB5AFD";
    when 16#085E# => romdata <= X"FAB0D701";
    when 16#085F# => romdata <= X"941DA548";
    when 16#0860# => romdata <= X"32FE8253";
    when 16#0861# => romdata <= X"BC0CF619";
    when 16#0862# => romdata <= X"24BCA2CA";
    when 16#0863# => romdata <= X"231A196C";
    when 16#0864# => romdata <= X"7C32A350";
    when 16#0865# => romdata <= X"AC9A5FA2";
    when 16#0866# => romdata <= X"884D8571";
    when 16#0867# => romdata <= X"FEEEDB7D";
    when 16#0868# => romdata <= X"29632E71";
    when 16#0869# => romdata <= X"898BB62B";
    when 16#086A# => romdata <= X"5E4E0104";
    when 16#086B# => romdata <= X"F73AA6A9";
    when 16#086C# => romdata <= X"C6B8CDA8";
    when 16#086D# => romdata <= X"16872805";
    when 16#086E# => romdata <= X"D75ECA64";
    when 16#086F# => romdata <= X"F9616410";
    when 16#0870# => romdata <= X"77B259C9";
    when 16#0871# => romdata <= X"D39E2F3C";
    when 16#0872# => romdata <= X"CD9FCFB1";
    when 16#0873# => romdata <= X"E6B6E269";
    when 16#0874# => romdata <= X"2EA34336";
    when 16#0875# => romdata <= X"A967E587";
    when 16#0876# => romdata <= X"F32E49B9";
    when 16#0877# => romdata <= X"61B91311";
    when 16#0878# => romdata <= X"198A204D";
    when 16#0879# => romdata <= X"11874B4B";
    when 16#087A# => romdata <= X"EBC6C04D";
    when 16#087B# => romdata <= X"DB5B82D5";
    when 16#087C# => romdata <= X"B741D3CE";
    when 16#087D# => romdata <= X"DC03A56A";
    when 16#087E# => romdata <= X"2017B3D2";
    when 16#087F# => romdata <= X"C4FBBD40";
    when 16#0880# => romdata <= X"CFDD6B78";
    when 16#0881# => romdata <= X"AEB21CDC";
    when 16#0882# => romdata <= X"D6AF8C34";
    when 16#0883# => romdata <= X"9F6DF8FF";
    when 16#0884# => romdata <= X"8B96BC82";
    when 16#0885# => romdata <= X"46A672A1";
    when 16#0886# => romdata <= X"6E45B5D0";
    when 16#0887# => romdata <= X"AB7D9925";
    when 16#0888# => romdata <= X"70EC45A5";
    when 16#0889# => romdata <= X"34B77F20";
    when 16#088A# => romdata <= X"4039FE20";
    when 16#088B# => romdata <= X"0D4C5E7C";
    when 16#088C# => romdata <= X"78FE2494";
    when 16#088D# => romdata <= X"1F578097";
    when 16#088E# => romdata <= X"B216177D";
    when 16#088F# => romdata <= X"8AD4E184";
    when 16#0890# => romdata <= X"4B2E52D8";
    when 16#0891# => romdata <= X"43256D0B";
    when 16#0892# => romdata <= X"E8504CF2";
    when 16#0893# => romdata <= X"D5B639E2";
    when 16#0894# => romdata <= X"CD501A6F";
    when 16#0895# => romdata <= X"E39B8AA7";
    when 16#0896# => romdata <= X"DB7DEA92";
    when 16#0897# => romdata <= X"4B38692E";
    when 16#0898# => romdata <= X"43195DB7";
    when 16#0899# => romdata <= X"E5F25E25";
    when 16#089A# => romdata <= X"152DF0FB";
    when 16#089B# => romdata <= X"7E0D4EF6";
    when 16#089C# => romdata <= X"3F99CD95";
    when 16#089D# => romdata <= X"F699E165";
    when 16#089E# => romdata <= X"76702B65";
    when 16#089F# => romdata <= X"1C295836";
    when 16#08A0# => romdata <= X"45070011";
    when 16#08A1# => romdata <= X"B2A1F88C";
    when 16#08A2# => romdata <= X"947BAE7C";
    when 16#08A3# => romdata <= X"94D48EB0";
    when 16#08A4# => romdata <= X"7A132DB3";
    when 16#08A5# => romdata <= X"8D4FE2B7";
    when 16#08A6# => romdata <= X"7EEAFB31";
    when 16#08A7# => romdata <= X"AFB44271";
    when 16#08A8# => romdata <= X"0BD0AE4E";
    when 16#08A9# => romdata <= X"6102DA69";
    when 16#08AA# => romdata <= X"A454517B";
    when 16#08AB# => romdata <= X"6F148D97";
    when 16#08AC# => romdata <= X"DBFBAC73";
    when 16#08AD# => romdata <= X"05979B5D";
    when 16#08AE# => romdata <= X"74D7D756";
    when 16#08AF# => romdata <= X"8A0CA56C";
    when 16#08B0# => romdata <= X"A89F23D8";
    when 16#08B1# => romdata <= X"33026102";
    when 16#08B2# => romdata <= X"5CC741F9";
    when 16#08B3# => romdata <= X"D7A4BDB3";
    when 16#08B4# => romdata <= X"56B544C6";
    when 16#08B5# => romdata <= X"8C89CCC2";
    when 16#08B6# => romdata <= X"C125F5C7";
    when 16#08B7# => romdata <= X"1E18C4EA";
    when 16#08B8# => romdata <= X"102343AE";
    when 16#08B9# => romdata <= X"4A44F6FC";
    when 16#08BA# => romdata <= X"695810E6";
    when 16#08BB# => romdata <= X"F28C86BF";
    when 16#08BC# => romdata <= X"53F4C8B8";
    when 16#08BD# => romdata <= X"AAE46DF6";
    when 16#08BE# => romdata <= X"006B1679";
    when 16#08BF# => romdata <= X"EBEA7902";
    when 16#08C0# => romdata <= X"66D4D02A";
    when 16#08C1# => romdata <= X"2095074A";
    when 16#08C2# => romdata <= X"DA634EE6";
    when 16#08C3# => romdata <= X"0C707028";
    when 16#08C4# => romdata <= X"5C316E1F";
    when 16#08C5# => romdata <= X"191BC5A8";
    when 16#08C6# => romdata <= X"8B80D673";
    when 16#08C7# => romdata <= X"F144D65B";
    when 16#08C8# => romdata <= X"870A65FC";
    when 16#08C9# => romdata <= X"93D8B4BB";
    when 16#08CA# => romdata <= X"29B80FD5";
    when 16#08CB# => romdata <= X"8F9FE95F";
    when 16#08CC# => romdata <= X"59948783";
    when 16#08CD# => romdata <= X"08CAC539";
    when 16#08CE# => romdata <= X"4781E4D5";
    when 16#08CF# => romdata <= X"A3F5EA2A";
    when 16#08D0# => romdata <= X"8ED834EE";
    when 16#08D1# => romdata <= X"5BD31D20";
    when 16#08D2# => romdata <= X"58C843F2";
    when 16#08D3# => romdata <= X"2EB778C4";
    when 16#08D4# => romdata <= X"C2514419";
    when 16#08D5# => romdata <= X"3DAA65F9";
    when 16#08D6# => romdata <= X"B57AEC4A";
    when 16#08D7# => romdata <= X"344713E9";
    when 16#08D8# => romdata <= X"EDF913F3";
    when 16#08D9# => romdata <= X"CD29196B";
    when 16#08DA# => romdata <= X"42E71BB1";
    when 16#08DB# => romdata <= X"82AC3B1A";
    when 16#08DC# => romdata <= X"60AFDBF1";
    when 16#08DD# => romdata <= X"112A86A2";
    when 16#08DE# => romdata <= X"0BFC1D28";
    when 16#08DF# => romdata <= X"D3E0DBBA";
    when 16#08E0# => romdata <= X"BF38E8F1";
    when 16#08E1# => romdata <= X"2651C207";
    when 16#08E2# => romdata <= X"C951654F";
    when 16#08E3# => romdata <= X"E8C4CECB";
    when 16#08E4# => romdata <= X"6C6F93EC";
    when 16#08E5# => romdata <= X"46456DAF";
    when 16#08E6# => romdata <= X"FD7320DE";
    when 16#08E7# => romdata <= X"C8D08F2F";
    when 16#08E8# => romdata <= X"712CEB4D";
    when 16#08E9# => romdata <= X"82407D61";
    when 16#08EA# => romdata <= X"CC47B333";
    when 16#08EB# => romdata <= X"F69310C0";
    when 16#08EC# => romdata <= X"6EE1FB5E";
    when 16#08ED# => romdata <= X"D84F8394";
    when 16#08EE# => romdata <= X"5F05D4A8";
    when 16#08EF# => romdata <= X"7CF5A68D";
    when 16#08F0# => romdata <= X"78B55368";
    when 16#08F1# => romdata <= X"80DE3443";
    when 16#08F2# => romdata <= X"E804040E";
    when 16#08F3# => romdata <= X"599BC583";
    when 16#08F4# => romdata <= X"7E22150C";
    when 16#08F5# => romdata <= X"93CC1E5E";
    when 16#08F6# => romdata <= X"711F9B88";
    when 16#08F7# => romdata <= X"9C78C6FF";
    when 16#08F8# => romdata <= X"882D8085";
    when 16#08F9# => romdata <= X"7EF41ABC";
    when 16#08FA# => romdata <= X"5F12E991";
    when 16#08FB# => romdata <= X"05E6C894";
    when 16#08FC# => romdata <= X"EC0B796E";
    when 16#08FD# => romdata <= X"0A645780";
    when 16#08FE# => romdata <= X"341CBD03";
    when 16#08FF# => romdata <= X"9E8C6EE0";
    when 16#0900# => romdata <= X"ABA759AE";
    when 16#0901# => romdata <= X"16B9D877";
    when 16#0902# => romdata <= X"8FAC203F";
    when 16#0903# => romdata <= X"ADF48015";
    when 16#0904# => romdata <= X"331D6499";
    when 16#0905# => romdata <= X"B8CD74BD";
    when 16#0906# => romdata <= X"71ABEBD3";
    when 16#0907# => romdata <= X"E53ED906";
    when 16#0908# => romdata <= X"25E3057E";
    when 16#0909# => romdata <= X"A47BE587";
    when 16#090A# => romdata <= X"600F308D";
    when 16#090B# => romdata <= X"38743A68";
    when 16#090C# => romdata <= X"6EF6FA18";
    when 16#090D# => romdata <= X"9A4D86E4";
    when 16#090E# => romdata <= X"A35EB798";
    when 16#090F# => romdata <= X"FD230734";
    when 16#0910# => romdata <= X"5FBD10FA";
    when 16#0911# => romdata <= X"701265F6";
    when 16#0912# => romdata <= X"41760336";
    when 16#0913# => romdata <= X"5FCC4CE7";
    when 16#0914# => romdata <= X"63592442";
    when 16#0915# => romdata <= X"8167115B";
    when 16#0916# => romdata <= X"A372294C";
    when 16#0917# => romdata <= X"27A23CE6";
    when 16#0918# => romdata <= X"C27C5066";
    when 16#0919# => romdata <= X"03C5A661";
    when 16#091A# => romdata <= X"8A2B3344";
    when 16#091B# => romdata <= X"BAC50AB7";
    when 16#091C# => romdata <= X"FDC29D36";
    when 16#091D# => romdata <= X"BCBDFCE0";
    when 16#091E# => romdata <= X"D48D088E";
    when 16#091F# => romdata <= X"FD8EA1DE";
    when 16#0920# => romdata <= X"492C5430";
    when 16#0921# => romdata <= X"93C30AB7";
    when 16#0922# => romdata <= X"694627C0";
    when 16#0923# => romdata <= X"1B334CE3";
    when 16#0924# => romdata <= X"368AEB4B";
    when 16#0925# => romdata <= X"B3267EBB";
    when 16#0926# => romdata <= X"1096450B";
    when 16#0927# => romdata <= X"DFC25719";
    when 16#0928# => romdata <= X"77D7EF78";
    when 16#0929# => romdata <= X"D6E288FC";
    when 16#092A# => romdata <= X"E0388A04";
    when 16#092B# => romdata <= X"1838EC20";
    when 16#092C# => romdata <= X"31248F5F";
    when 16#092D# => romdata <= X"D659C701";
    when 16#092E# => romdata <= X"80634A1D";
    when 16#092F# => romdata <= X"C7196C8D";
    when 16#0930# => romdata <= X"9111C75B";
    when 16#0931# => romdata <= X"51C50F85";
    when 16#0932# => romdata <= X"4CEC63DE";
    when 16#0933# => romdata <= X"BF9FFE1A";
    when 16#0934# => romdata <= X"B9406735";
    when 16#0935# => romdata <= X"EC318727";
    when 16#0936# => romdata <= X"6DE7CA2F";
    when 16#0937# => romdata <= X"AD428702";
    when 16#0938# => romdata <= X"7956C93B";
    when 16#0939# => romdata <= X"8E84B7C0";
    when 16#093A# => romdata <= X"C3A9C3F7";
    when 16#093B# => romdata <= X"E82B3DB3";
    when 16#093C# => romdata <= X"5EB6D2CE";
    when 16#093D# => romdata <= X"BDFE0708";
    when 16#093E# => romdata <= X"FEDD764C";
    when 16#093F# => romdata <= X"839954F2";
    when 16#0940# => romdata <= X"CC9044B6";
    when 16#0941# => romdata <= X"52D0A01D";
    when 16#0942# => romdata <= X"28BD6B9D";
    when 16#0943# => romdata <= X"3DD9740C";
    when 16#0944# => romdata <= X"AE39AA52";
    when 16#0945# => romdata <= X"597FFC12";
    when 16#0946# => romdata <= X"27FAD8B7";
    when 16#0947# => romdata <= X"8EAFFC31";
    when 16#0948# => romdata <= X"BE94A632";
    when 16#0949# => romdata <= X"A1AA7A60";
    when 16#094A# => romdata <= X"AA5A9E09";
    when 16#094B# => romdata <= X"0DA2B62F";
    when 16#094C# => romdata <= X"6DBDFDC5";
    when 16#094D# => romdata <= X"0DF6EBE1";
    when 16#094E# => romdata <= X"D9949619";
    when 16#094F# => romdata <= X"FE9B2302";
    when 16#0950# => romdata <= X"248D6C80";
    when 16#0951# => romdata <= X"1DD2D6C0";
    when 16#0952# => romdata <= X"1FF8206A";
    when 16#0953# => romdata <= X"93C0AD22";
    when 16#0954# => romdata <= X"C6990C4E";
    when 16#0955# => romdata <= X"ECA7D4BD";
    when 16#0956# => romdata <= X"F36C3246";
    when 16#0957# => romdata <= X"A5D2D2B3";
    when 16#0958# => romdata <= X"982C608E";
    when 16#0959# => romdata <= X"6AD6BDD8";
    when 16#095A# => romdata <= X"5C92682E";
    when 16#095B# => romdata <= X"BDC9E411";
    when 16#095C# => romdata <= X"7F8B7F84";
    when 16#095D# => romdata <= X"1239C2A5";
    when 16#095E# => romdata <= X"AD7977E1";
    when 16#095F# => romdata <= X"1E4E9CA7";
    when 16#0960# => romdata <= X"3A55859E";
    when 16#0961# => romdata <= X"ADF7C9C2";
    when 16#0962# => romdata <= X"F1B28A6B";
    when 16#0963# => romdata <= X"4AC72020";
    when 16#0964# => romdata <= X"19230063";
    when 16#0965# => romdata <= X"331FC558";
    when 16#0966# => romdata <= X"6756CEA1";
    when 16#0967# => romdata <= X"F8478173";
    when 16#0968# => romdata <= X"A0A4964D";
    when 16#0969# => romdata <= X"00C1AC09";
    when 16#096A# => romdata <= X"95901521";
    when 16#096B# => romdata <= X"25A4D015";
    when 16#096C# => romdata <= X"92C54DC2";
    when 16#096D# => romdata <= X"555E1BA3";
    when 16#096E# => romdata <= X"4C7AC039";
    when 16#096F# => romdata <= X"394D1979";
    when 16#0970# => romdata <= X"AEA2BF7B";
    when 16#0971# => romdata <= X"2B2A8CB9";
    when 16#0972# => romdata <= X"D62E8913";
    when 16#0973# => romdata <= X"2CE9E3B3";
    when 16#0974# => romdata <= X"25F023AC";
    when 16#0975# => romdata <= X"6E8117CE";
    when 16#0976# => romdata <= X"57AD4B27";
    when 16#0977# => romdata <= X"1EFB0C17";
    when 16#0978# => romdata <= X"2FBFF8FA";
    when 16#0979# => romdata <= X"6A17A490";
    when 16#097A# => romdata <= X"B67CA7B1";
    when 16#097B# => romdata <= X"5F865A8A";
    when 16#097C# => romdata <= X"EEF37651";
    when 16#097D# => romdata <= X"A622390E";
    when 16#097E# => romdata <= X"82AFD418";
    when 16#097F# => romdata <= X"C7AFD480";
    when 16#0980# => romdata <= X"CEA29601";
    when 16#0981# => romdata <= X"B96AD3A8";
    when 16#0982# => romdata <= X"31646922";
    when 16#0983# => romdata <= X"000BBFF0";
    when 16#0984# => romdata <= X"2C014A91";
    when 16#0985# => romdata <= X"36D9A151";
    when 16#0986# => romdata <= X"A0E61A51";
    when 16#0987# => romdata <= X"F9FC2EC0";
    when 16#0988# => romdata <= X"C3A8F4C8";
    when 16#0989# => romdata <= X"3E64BDE5";
    when 16#098A# => romdata <= X"69A33B4C";
    when 16#098B# => romdata <= X"D653C134";
    when 16#098C# => romdata <= X"5B7CBEA3";
    when 16#098D# => romdata <= X"B3AC0411";
    when 16#098E# => romdata <= X"B6145727";
    when 16#098F# => romdata <= X"B1DBF606";
    when 16#0990# => romdata <= X"6ABCE9DA";
    when 16#0991# => romdata <= X"A8B0DE58";
    when 16#0992# => romdata <= X"ADC2510C";
    when 16#0993# => romdata <= X"02C2619A";
    when 16#0994# => romdata <= X"542A139F";
    when 16#0995# => romdata <= X"A3EF7A03";
    when 16#0996# => romdata <= X"AD346734";
    when 16#0997# => romdata <= X"5D9573C1";
    when 16#0998# => romdata <= X"07A13E7F";
    when 16#0999# => romdata <= X"CD43C0D5";
    when 16#099A# => romdata <= X"1DB5EC1A";
    when 16#099B# => romdata <= X"09D409DA";
    when 16#099C# => romdata <= X"75462F9C";
    when 16#099D# => romdata <= X"71F0C9E3";
    when 16#099E# => romdata <= X"6C2742C2";
    when 16#099F# => romdata <= X"79C910F0";
    when 16#09A0# => romdata <= X"7CFC5CF7";
    when 16#09A1# => romdata <= X"F98AD48D";
    when 16#09A2# => romdata <= X"67232A2D";
    when 16#09A3# => romdata <= X"F29A66B7";
    when 16#09A4# => romdata <= X"82095573";
    when 16#09A5# => romdata <= X"57A4BC91";
    when 16#09A6# => romdata <= X"922D4195";
    when 16#09A7# => romdata <= X"DA9533CD";
    when 16#09A8# => romdata <= X"3501F388";
    when 16#09A9# => romdata <= X"AF6EE2BB";
    when 16#09AA# => romdata <= X"3AD08BC7";
    when 16#09AB# => romdata <= X"D5301505";
    when 16#09AC# => romdata <= X"9988F5B9";
    when 16#09AD# => romdata <= X"BF7824D0";
    when 16#09AE# => romdata <= X"66DCBDC6";
    when 16#09AF# => romdata <= X"1CA588DC";
    when 16#09B0# => romdata <= X"CF0EBDE4";
    when 16#09B1# => romdata <= X"A96632DB";
    when 16#09B2# => romdata <= X"A22CA0D7";
    when 16#09B3# => romdata <= X"70C61A1D";
    when 16#09B4# => romdata <= X"D66EDA88";
    when 16#09B5# => romdata <= X"2D02C5FA";
    when 16#09B6# => romdata <= X"284798E1";
    when 16#09B7# => romdata <= X"2296E89C";
    when 16#09B8# => romdata <= X"45906D31";
    when 16#09B9# => romdata <= X"5EFDBA81";
    when 16#09BA# => romdata <= X"6FD869DF";
    when 16#09BB# => romdata <= X"869A65DD";
    when 16#09BC# => romdata <= X"8BA4E0B1";
    when 16#09BD# => romdata <= X"3C441EEB";
    when 16#09BE# => romdata <= X"052EF3D0";
    when 16#09BF# => romdata <= X"FD436E4A";
    when 16#09C0# => romdata <= X"C68EFC74";
    when 16#09C1# => romdata <= X"9E0CF4C7";
    when 16#09C2# => romdata <= X"E15599D5";
    when 16#09C3# => romdata <= X"514E136A";
    when 16#09C4# => romdata <= X"BD134BA6";
    when 16#09C5# => romdata <= X"38A02E9E";
    when 16#09C6# => romdata <= X"C1FE66CC";
    when 16#09C7# => romdata <= X"9ACBCE50";
    when 16#09C8# => romdata <= X"82C87341";
    when 16#09C9# => romdata <= X"96BADC21";
    when 16#09CA# => romdata <= X"F4DA7621";
    when 16#09CB# => romdata <= X"D9FA7253";
    when 16#09CC# => romdata <= X"62C41112";
    when 16#09CD# => romdata <= X"7836A26C";
    when 16#09CE# => romdata <= X"B44CB385";
    when 16#09CF# => romdata <= X"1D53C599";
    when 16#09D0# => romdata <= X"B94A5E67";
    when 16#09D1# => romdata <= X"862665D7";
    when 16#09D2# => romdata <= X"092C43D9";
    when 16#09D3# => romdata <= X"B4AD3FE2";
    when 16#09D4# => romdata <= X"0B8AFACC";
    when 16#09D5# => romdata <= X"EDE920F4";
    when 16#09D6# => romdata <= X"40F3BF55";
    when 16#09D7# => romdata <= X"52CFAFAD";
    when 16#09D8# => romdata <= X"04A7D7E0";
    when 16#09D9# => romdata <= X"A9CEA18D";
    when 16#09DA# => romdata <= X"497282D4";
    when 16#09DB# => romdata <= X"4778FB7D";
    when 16#09DC# => romdata <= X"5072832C";
    when 16#09DD# => romdata <= X"0B77C4C5";
    when 16#09DE# => romdata <= X"1F4DCFD7";
    when 16#09DF# => romdata <= X"AC07DC7A";
    when 16#09E0# => romdata <= X"9863DB8A";
    when 16#09E1# => romdata <= X"38F1C003";
    when 16#09E2# => romdata <= X"CB852F61";
    when 16#09E3# => romdata <= X"19BE801A";
    when 16#09E4# => romdata <= X"D12B8BC7";
    when 16#09E5# => romdata <= X"393B0064";
    when 16#09E6# => romdata <= X"0F125C73";
    when 16#09E7# => romdata <= X"4447DB2F";
    when 16#09E8# => romdata <= X"D8B02F7F";
    when 16#09E9# => romdata <= X"7FC7A23B";
    when 16#09EA# => romdata <= X"84FB80F9";
    when 16#09EB# => romdata <= X"CC08E3EF";
    when 16#09EC# => romdata <= X"888634FF";
    when 16#09ED# => romdata <= X"B6F51ECE";
    when 16#09EE# => romdata <= X"E9B20A89";
    when 16#09EF# => romdata <= X"941FBF2B";
    when 16#09F0# => romdata <= X"49314DBD";
    when 16#09F1# => romdata <= X"D67CB7A1";
    when 16#09F2# => romdata <= X"B5BD8D62";
    when 16#09F3# => romdata <= X"9FA327AF";
    when 16#09F4# => romdata <= X"2CBB47B5";
    when 16#09F5# => romdata <= X"419A0A8C";
    when 16#09F6# => romdata <= X"B807D301";
    when 16#09F7# => romdata <= X"52FA5606";
    when 16#09F8# => romdata <= X"90DBAC49";
    when 16#09F9# => romdata <= X"D6B043D5";
    when 16#09FA# => romdata <= X"BC9D51E8";
    when 16#09FB# => romdata <= X"2C3B1CF4";
    when 16#09FC# => romdata <= X"ED69E997";
    when 16#09FD# => romdata <= X"050C6519";
    when 16#09FE# => romdata <= X"7F3D93E2";
    when 16#09FF# => romdata <= X"1CBE91E0";
    when 16#0A00# => romdata <= X"D358BFC8";
    when 16#0A01# => romdata <= X"C6AD1DC9";
    when 16#0A02# => romdata <= X"4E71D1F5";
    when 16#0A03# => romdata <= X"D0558942";
    when 16#0A04# => romdata <= X"4275875A";
    when 16#0A05# => romdata <= X"F8CDA2AB";
    when 16#0A06# => romdata <= X"CC6404D6";
    when 16#0A07# => romdata <= X"FCB7A2E0";
    when 16#0A08# => romdata <= X"A74C6802";
    when 16#0A09# => romdata <= X"4827E026";
    when 16#0A0A# => romdata <= X"21C10CD5";
    when 16#0A0B# => romdata <= X"FB149FBA";
    when 16#0A0C# => romdata <= X"373AE32D";
    when 16#0A0D# => romdata <= X"FFF275CF";
    when 16#0A0E# => romdata <= X"386C3D7A";
    when 16#0A0F# => romdata <= X"04E3FE10";
    when 16#0A10# => romdata <= X"B6F1A6F4";
    when 16#0A11# => romdata <= X"782B4823";
    when 16#0A12# => romdata <= X"242F2967";
    when 16#0A13# => romdata <= X"2E847CCE";
    when 16#0A14# => romdata <= X"760BA005";
    when 16#0A15# => romdata <= X"D6852A34";
    when 16#0A16# => romdata <= X"59E7576A";
    when 16#0A17# => romdata <= X"254B10A9";
    when 16#0A18# => romdata <= X"A78A9F81";
    when 16#0A19# => romdata <= X"12BEA39B";
    when 16#0A1A# => romdata <= X"A65898CF";
    when 16#0A1B# => romdata <= X"ED1179D6";
    when 16#0A1C# => romdata <= X"8211D98E";
    when 16#0A1D# => romdata <= X"6950ED06";
    when 16#0A1E# => romdata <= X"399E3943";
    when 16#0A1F# => romdata <= X"3ACD898E";
    when 16#0A20# => romdata <= X"2F6C87F5";
    when 16#0A21# => romdata <= X"FB9D9951";
    when 16#0A22# => romdata <= X"8EF36429";
    when 16#0A23# => romdata <= X"D447B0EF";
    when 16#0A24# => romdata <= X"0C5B7D83";
    when 16#0A25# => romdata <= X"4ACFA388";
    when 16#0A26# => romdata <= X"578BDF60";
    when 16#0A27# => romdata <= X"D4B1FB5A";
    when 16#0A28# => romdata <= X"0CEE7D1D";
    when 16#0A29# => romdata <= X"613BB9B9";
    when 16#0A2A# => romdata <= X"9E36DC96";
    when 16#0A2B# => romdata <= X"36E70A54";
    when 16#0A2C# => romdata <= X"3BA6BF0B";
    when 16#0A2D# => romdata <= X"3A448DBD";
    when 16#0A2E# => romdata <= X"F8046949";
    when 16#0A2F# => romdata <= X"4239D4B7";
    when 16#0A30# => romdata <= X"C4979D82";
    when 16#0A31# => romdata <= X"E80C08EF";
    when 16#0A32# => romdata <= X"36EA6756";
    when 16#0A33# => romdata <= X"0C86665D";
    when 16#0A34# => romdata <= X"458040CE";
    when 16#0A35# => romdata <= X"31BA009B";
    when 16#0A36# => romdata <= X"CDC30CCB";
    when 16#0A37# => romdata <= X"AC50259E";
    when 16#0A38# => romdata <= X"4485E570";
    when 16#0A39# => romdata <= X"F190613C";
    when 16#0A3A# => romdata <= X"B010563F";
    when 16#0A3B# => romdata <= X"6BD24C2F";
    when 16#0A3C# => romdata <= X"1CF73F6A";
    when 16#0A3D# => romdata <= X"6844AB83";
    when 16#0A3E# => romdata <= X"50D23BBC";
    when 16#0A3F# => romdata <= X"3D1361E7";
    when 16#0A40# => romdata <= X"3DCE94AF";
    when 16#0A41# => romdata <= X"83697BB8";
    when 16#0A42# => romdata <= X"17BA366C";
    when 16#0A43# => romdata <= X"9855A754";
    when 16#0A44# => romdata <= X"EFC2F007";
    when 16#0A45# => romdata <= X"D99A9641";
    when 16#0A46# => romdata <= X"25682E6F";
    when 16#0A47# => romdata <= X"5CF7FBBF";
    when 16#0A48# => romdata <= X"687D221B";
    when 16#0A49# => romdata <= X"5A0FD844";
    when 16#0A4A# => romdata <= X"477A2F87";
    when 16#0A4B# => romdata <= X"D5370F44";
    when 16#0A4C# => romdata <= X"69F76073";
    when 16#0A4D# => romdata <= X"A93AEF78";
    when 16#0A4E# => romdata <= X"12275FD4";
    when 16#0A4F# => romdata <= X"F70B2040";
    when 16#0A50# => romdata <= X"C12A83AD";
    when 16#0A51# => romdata <= X"E5E5D862";
    when 16#0A52# => romdata <= X"684D119D";
    when 16#0A53# => romdata <= X"CA0F75AE";
    when 16#0A54# => romdata <= X"2B56C794";
    when 16#0A55# => romdata <= X"968A6856";
    when 16#0A56# => romdata <= X"6291B731";
    when 16#0A57# => romdata <= X"579A1055";
    when 16#0A58# => romdata <= X"A84F083B";
    when 16#0A59# => romdata <= X"3072B7BD";
    when 16#0A5A# => romdata <= X"5AC9D520";
    when 16#0A5B# => romdata <= X"F64F0829";
    when 16#0A5C# => romdata <= X"B5928756";
    when 16#0A5D# => romdata <= X"13BDD81C";
    when 16#0A5E# => romdata <= X"11622B33";
    when 16#0A5F# => romdata <= X"1289C985";
    when 16#0A60# => romdata <= X"01B01EE1";
    when 16#0A61# => romdata <= X"D813C0E9";
    when 16#0A62# => romdata <= X"7CF36878";
    when 16#0A63# => romdata <= X"260F80BF";
    when 16#0A64# => romdata <= X"88071D25";
    when 16#0A65# => romdata <= X"8B9DE02F";
    when 16#0A66# => romdata <= X"3F90B4C1";
    when 16#0A67# => romdata <= X"2BB56CBC";
    when 16#0A68# => romdata <= X"731550B5";
    when 16#0A69# => romdata <= X"EFDE6D97";
    when 16#0A6A# => romdata <= X"A1283EEF";
    when 16#0A6B# => romdata <= X"E61CD6E5";
    when 16#0A6C# => romdata <= X"DF312D0F";
    when 16#0A6D# => romdata <= X"0153A32D";
    when 16#0A6E# => romdata <= X"D65B143E";
    when 16#0A6F# => romdata <= X"C6A3F2B6";
    when 16#0A70# => romdata <= X"4E2B8FFB";
    when 16#0A71# => romdata <= X"47EAE46B";
    when 16#0A72# => romdata <= X"D92A6EB9";
    when 16#0A73# => romdata <= X"ACBDD11A";
    when 16#0A74# => romdata <= X"2D730D02";
    when 16#0A75# => romdata <= X"7A3EDEAD";
    when 16#0A76# => romdata <= X"BA596519";
    when 16#0A77# => romdata <= X"8FD59BBC";
    when 16#0A78# => romdata <= X"8574B680";
    when 16#0A79# => romdata <= X"B96AD485";
    when 16#0A7A# => romdata <= X"86E5B176";
    when 16#0A7B# => romdata <= X"25251BF4";
    when 16#0A7C# => romdata <= X"374E28C6";
    when 16#0A7D# => romdata <= X"AB956C68";
    when 16#0A7E# => romdata <= X"18183FDC";
    when 16#0A7F# => romdata <= X"119499E0";
    when 16#0A80# => romdata <= X"FE694332";
    when 16#0A81# => romdata <= X"33B6067B";
    when 16#0A82# => romdata <= X"0EACF1F4";
    when 16#0A83# => romdata <= X"7BD3AAD9";
    when 16#0A84# => romdata <= X"783FA30F";
    when 16#0A85# => romdata <= X"684110D1";
    when 16#0A86# => romdata <= X"15245923";
    when 16#0A87# => romdata <= X"3896479D";
    when 16#0A88# => romdata <= X"08A976B8";
    when 16#0A89# => romdata <= X"53E4B7B5";
    when 16#0A8A# => romdata <= X"2A345112";
    when 16#0A8B# => romdata <= X"39961048";
    when 16#0A8C# => romdata <= X"B7C1B900";
    when 16#0A8D# => romdata <= X"9095327C";
    when 16#0A8E# => romdata <= X"86F2EA29";
    when 16#0A8F# => romdata <= X"1FAC1734";
    when 16#0A90# => romdata <= X"ED2596EF";
    when 16#0A91# => romdata <= X"19D04528";
    when 16#0A92# => romdata <= X"F3D8F2A3";
    when 16#0A93# => romdata <= X"430A0C19";
    when 16#0A94# => romdata <= X"DA6A70A3";
    when 16#0A95# => romdata <= X"7DB6DC03";
    when 16#0A96# => romdata <= X"4BA0053B";
    when 16#0A97# => romdata <= X"57ACB9E7";
    when 16#0A98# => romdata <= X"C00ED9BD";
    when 16#0A99# => romdata <= X"6AC11339";
    when 16#0A9A# => romdata <= X"EA169D9D";
    when 16#0A9B# => romdata <= X"54E6739B";
    when 16#0A9C# => romdata <= X"051AF40E";
    when 16#0A9D# => romdata <= X"E79A1034";
    when 16#0A9E# => romdata <= X"D6294261";
    when 16#0A9F# => romdata <= X"E1AFFCD6";
    when 16#0AA0# => romdata <= X"1B9CA501";
    when 16#0AA1# => romdata <= X"6C56B2D1";
    when 16#0AA2# => romdata <= X"172D9B2A";
    when 16#0AA3# => romdata <= X"7283E4EE";
    when 16#0AA4# => romdata <= X"0A06C814";
    when 16#0AA5# => romdata <= X"9E5A2DAA";
    when 16#0AA6# => romdata <= X"263A5D24";
    when 16#0AA7# => romdata <= X"29C2B1FC";
    when 16#0AA8# => romdata <= X"E75C4188";
    when 16#0AA9# => romdata <= X"7DD02E05";
    when 16#0AAA# => romdata <= X"6EF87246";
    when 16#0AAB# => romdata <= X"45FEC6FE";
    when 16#0AAC# => romdata <= X"7FC1EF18";
    when 16#0AAD# => romdata <= X"0529B1E8";
    when 16#0AAE# => romdata <= X"94773CF3";
    when 16#0AAF# => romdata <= X"E2E1D938";
    when 16#0AB0# => romdata <= X"EFE9CD82";
    when 16#0AB1# => romdata <= X"4D914541";
    when 16#0AB2# => romdata <= X"16797F5A";
    when 16#0AB3# => romdata <= X"84746537";
    when 16#0AB4# => romdata <= X"FED5F0EB";
    when 16#0AB5# => romdata <= X"F0583C85";
    when 16#0AB6# => romdata <= X"08EA0745";
    when 16#0AB7# => romdata <= X"B4989954";
    when 16#0AB8# => romdata <= X"EBC4F215";
    when 16#0AB9# => romdata <= X"BE3D5156";
    when 16#0ABA# => romdata <= X"87BCDD5D";
    when 16#0ABB# => romdata <= X"FDAB9814";
    when 16#0ABC# => romdata <= X"358B0703";
    when 16#0ABD# => romdata <= X"8E0CB869";
    when 16#0ABE# => romdata <= X"A8C34F91";
    when 16#0ABF# => romdata <= X"6FC67773";
    when 16#0AC0# => romdata <= X"191679C6";
    when 16#0AC1# => romdata <= X"0A15A0A3";
    when 16#0AC2# => romdata <= X"99E224D0";
    when 16#0AC3# => romdata <= X"B0168439";
    when 16#0AC4# => romdata <= X"386C0AEE";
    when 16#0AC5# => romdata <= X"8F5EF771";
    when 16#0AC6# => romdata <= X"85AC847A";
    when 16#0AC7# => romdata <= X"66D934CB";
    when 16#0AC8# => romdata <= X"0ED6A346";
    when 16#0AC9# => romdata <= X"7C3B386B";
    when 16#0ACA# => romdata <= X"A7F11587";
    when 16#0ACB# => romdata <= X"7F36B49E";
    when 16#0ACC# => romdata <= X"111DE49E";
    when 16#0ACD# => romdata <= X"409468F3";
    when 16#0ACE# => romdata <= X"43A98974";
    when 16#0ACF# => romdata <= X"F4EF1EEE";
    when 16#0AD0# => romdata <= X"DD282F73";
    when 16#0AD1# => romdata <= X"013EC272";
    when 16#0AD2# => romdata <= X"7518DB46";
    when 16#0AD3# => romdata <= X"C6751A58";
    when 16#0AD4# => romdata <= X"AE3E0D5F";
    when 16#0AD5# => romdata <= X"9D2B966D";
    when 16#0AD6# => romdata <= X"4465BC55";
    when 16#0AD7# => romdata <= X"95BC31B2";
    when 16#0AD8# => romdata <= X"712AE1E1";
    when 16#0AD9# => romdata <= X"BF9915CC";
    when 16#0ADA# => romdata <= X"0E02CA72";
    when 16#0ADB# => romdata <= X"40EBB9A0";
    when 16#0ADC# => romdata <= X"45F959E7";
    when 16#0ADD# => romdata <= X"7DFCDADA";
    when 16#0ADE# => romdata <= X"B6248D58";
    when 16#0ADF# => romdata <= X"B47BBEF3";
    when 16#0AE0# => romdata <= X"C775DEFD";
    when 16#0AE1# => romdata <= X"629A2EED";
    when 16#0AE2# => romdata <= X"15201A21";
    when 16#0AE3# => romdata <= X"ADCA470B";
    when 16#0AE4# => romdata <= X"1AD30849";
    when 16#0AE5# => romdata <= X"24FABCDA";
    when 16#0AE6# => romdata <= X"B6B12FA6";
    when 16#0AE7# => romdata <= X"201E2A23";
    when 16#0AE8# => romdata <= X"9AE8F1BC";
    when 16#0AE9# => romdata <= X"D7CC39FE";
    when 16#0AEA# => romdata <= X"C62587E5";
    when 16#0AEB# => romdata <= X"8C84AAC1";
    when 16#0AEC# => romdata <= X"5935D452";
    when 16#0AED# => romdata <= X"61E3AFEB";
    when 16#0AEE# => romdata <= X"60016AFA";
    when 16#0AEF# => romdata <= X"0902DB98";
    when 16#0AF0# => romdata <= X"DCFE5865";
    when 16#0AF1# => romdata <= X"13FF70EF";
    when 16#0AF2# => romdata <= X"4E3F4777";
    when 16#0AF3# => romdata <= X"3635D475";
    when 16#0AF4# => romdata <= X"754A158F";
    when 16#0AF5# => romdata <= X"ACC9C470";
    when 16#0AF6# => romdata <= X"921FB018";
    when 16#0AF7# => romdata <= X"6BD6EEDE";
    when 16#0AF8# => romdata <= X"FCBEE9C8";
    when 16#0AF9# => romdata <= X"03118851";
    when 16#0AFA# => romdata <= X"F82CACBF";
    when 16#0AFB# => romdata <= X"8C0A544B";
    when 16#0AFC# => romdata <= X"0562E2E2";
    when 16#0AFD# => romdata <= X"7286CEA5";
    when 16#0AFE# => romdata <= X"FBAF83AA";
    when 16#0AFF# => romdata <= X"5C1F97A0";
    when 16#0B00# => romdata <= X"C7386F9F";
    when 16#0B01# => romdata <= X"F39FDDBF";
    when 16#0B02# => romdata <= X"EB223AD8";
    when 16#0B03# => romdata <= X"B856EA2E";
    when 16#0B04# => romdata <= X"7F3AFEDE";
    when 16#0B05# => romdata <= X"197A61F1";
    when 16#0B06# => romdata <= X"83FF7DF2";
    when 16#0B07# => romdata <= X"FD6DE208";
    when 16#0B08# => romdata <= X"E71E6E10";
    when 16#0B09# => romdata <= X"63FB3774";
    when 16#0B0A# => romdata <= X"B6969135";
    when 16#0B0B# => romdata <= X"24F7488E";
    when 16#0B0C# => romdata <= X"FC2CA54E";
    when 16#0B0D# => romdata <= X"8B653EF5";
    when 16#0B0E# => romdata <= X"BCB7A8F4";
    when 16#0B0F# => romdata <= X"994E312D";
    when 16#0B10# => romdata <= X"CEE99A31";
    when 16#0B11# => romdata <= X"6C2ABF3F";
    when 16#0B12# => romdata <= X"DF85B8FA";
    when 16#0B13# => romdata <= X"9BBD4366";
    when 16#0B14# => romdata <= X"ABBD7B3D";
    when 16#0B15# => romdata <= X"3D433C14";
    when 16#0B16# => romdata <= X"710A95EB";
    when 16#0B17# => romdata <= X"B3D0FCDA";
    when 16#0B18# => romdata <= X"2D37A443";
    when 16#0B19# => romdata <= X"D62A8361";
    when 16#0B1A# => romdata <= X"DA78ACA7";
    when 16#0B1B# => romdata <= X"81CEC045";
    when 16#0B1C# => romdata <= X"42D01DE7";
    when 16#0B1D# => romdata <= X"B6C6D14C";
    when 16#0B1E# => romdata <= X"DD4EA709";
    when 16#0B1F# => romdata <= X"264251D4";
    when 16#0B20# => romdata <= X"6C42AAF4";
    when 16#0B21# => romdata <= X"04094286";
    when 16#0B22# => romdata <= X"DA5BFF8E";
    when 16#0B23# => romdata <= X"81FA2F8C";
    when 16#0B24# => romdata <= X"54B17282";
    when 16#0B25# => romdata <= X"1054F4CE";
    when 16#0B26# => romdata <= X"D82287F2";
    when 16#0B27# => romdata <= X"9EA3D3AA";
    when 16#0B28# => romdata <= X"798C9CF5";
    when 16#0B29# => romdata <= X"C5A909B9";
    when 16#0B2A# => romdata <= X"FBA641A8";
    when 16#0B2B# => romdata <= X"D9E31024";
    when 16#0B2C# => romdata <= X"8B0F9A13";
    when 16#0B2D# => romdata <= X"75CE4DAA";
    when 16#0B2E# => romdata <= X"98EB6228";
    when 16#0B2F# => romdata <= X"6B4EF4DF";
    when 16#0B30# => romdata <= X"C58B877A";
    when 16#0B31# => romdata <= X"73D017B1";
    when 16#0B32# => romdata <= X"7AFD7F1F";
    when 16#0B33# => romdata <= X"58D3D2CA";
    when 16#0B34# => romdata <= X"D3B7AF2F";
    when 16#0B35# => romdata <= X"06699B08";
    when 16#0B36# => romdata <= X"B88FB4EB";
    when 16#0B37# => romdata <= X"70D25111";
    when 16#0B38# => romdata <= X"90158BB4";
    when 16#0B39# => romdata <= X"928ED173";
    when 16#0B3A# => romdata <= X"5C944009";
    when 16#0B3B# => romdata <= X"80144EF9";
    when 16#0B3C# => romdata <= X"ED06E060";
    when 16#0B3D# => romdata <= X"74E2F293";
    when 16#0B3E# => romdata <= X"25C1AA31";
    when 16#0B3F# => romdata <= X"6A46E8E6";
    when 16#0B40# => romdata <= X"17B3CE91";
    when 16#0B41# => romdata <= X"6CFCF05A";
    when 16#0B42# => romdata <= X"389052DE";
    when 16#0B43# => romdata <= X"12049834";
    when 16#0B44# => romdata <= X"1EE26A27";
    when 16#0B45# => romdata <= X"A3D757AA";
    when 16#0B46# => romdata <= X"E763046B";
    when 16#0B47# => romdata <= X"8CBC8413";
    when 16#0B48# => romdata <= X"50292F06";
    when 16#0B49# => romdata <= X"AFF97C97";
    when 16#0B4A# => romdata <= X"07CE5561";
    when 16#0B4B# => romdata <= X"F5C119E2";
    when 16#0B4C# => romdata <= X"FF6C1370";
    when 16#0B4D# => romdata <= X"94F62573";
    when 16#0B4E# => romdata <= X"EB80DC13";
    when 16#0B4F# => romdata <= X"862797C3";
    when 16#0B50# => romdata <= X"319158DD";
    when 16#0B51# => romdata <= X"D465FBC0";
    when 16#0B52# => romdata <= X"33CAD81B";
    when 16#0B53# => romdata <= X"FBBBB54D";
    when 16#0B54# => romdata <= X"9467599D";
    when 16#0B55# => romdata <= X"751B9980";
    when 16#0B56# => romdata <= X"A9AE8BFC";
    when 16#0B57# => romdata <= X"6715C5EA";
    when 16#0B58# => romdata <= X"74859E6A";
    when 16#0B59# => romdata <= X"10DB369D";
    when 16#0B5A# => romdata <= X"5DF83A92";
    when 16#0B5B# => romdata <= X"655A9A59";
    when 16#0B5C# => romdata <= X"08228B33";
    when 16#0B5D# => romdata <= X"B36F55DE";
    when 16#0B5E# => romdata <= X"563005B8";
    when 16#0B5F# => romdata <= X"86EB324C";
    when 16#0B60# => romdata <= X"EC4160F0";
    when 16#0B61# => romdata <= X"D18938E9";
    when 16#0B62# => romdata <= X"FE41D392";
    when 16#0B63# => romdata <= X"34C29E13";
    when 16#0B64# => romdata <= X"B814DDCD";
    when 16#0B65# => romdata <= X"13CA6450";
    when 16#0B66# => romdata <= X"77480092";
    when 16#0B67# => romdata <= X"4B084873";
    when 16#0B68# => romdata <= X"5C5DE076";
    when 16#0B69# => romdata <= X"F66EDC97";
    when 16#0B6A# => romdata <= X"3FC83B13";
    when 16#0B6B# => romdata <= X"938811CD";
    when 16#0B6C# => romdata <= X"98873714";
    when 16#0B6D# => romdata <= X"70AC5DD9";
    when 16#0B6E# => romdata <= X"85481185";
    when 16#0B6F# => romdata <= X"F1191EA8";
    when 16#0B70# => romdata <= X"C1D3A7DC";
    when 16#0B71# => romdata <= X"65E1E82E";
    when 16#0B72# => romdata <= X"2318D0FF";
    when 16#0B73# => romdata <= X"0C9AF65E";
    when 16#0B74# => romdata <= X"A1515DDC";
    when 16#0B75# => romdata <= X"536C5A8B";
    when 16#0B76# => romdata <= X"D0AF4817";
    when 16#0B77# => romdata <= X"89838DA5";
    when 16#0B78# => romdata <= X"4A39BA56";
    when 16#0B79# => romdata <= X"D014E122";
    when 16#0B7A# => romdata <= X"42600AC7";
    when 16#0B7B# => romdata <= X"8D28ADAC";
    when 16#0B7C# => romdata <= X"3FFD3600";
    when 16#0B7D# => romdata <= X"E8964458";
    when 16#0B7E# => romdata <= X"68064D1D";
    when 16#0B7F# => romdata <= X"2ACF22E0";
    when 16#0B80# => romdata <= X"BF5202D3";
    when 16#0B81# => romdata <= X"599D2DDA";
    when 16#0B82# => romdata <= X"AE5F526B";
    when 16#0B83# => romdata <= X"6B6AC469";
    when 16#0B84# => romdata <= X"D4BA0D0B";
    when 16#0B85# => romdata <= X"A5D79B1D";
    when 16#0B86# => romdata <= X"B8917332";
    when 16#0B87# => romdata <= X"0F0EB68F";
    when 16#0B88# => romdata <= X"5D9DA495";
    when 16#0B89# => romdata <= X"AA0981F8";
    when 16#0B8A# => romdata <= X"022426F6";
    when 16#0B8B# => romdata <= X"8519B548";
    when 16#0B8C# => romdata <= X"B19B5F8C";
    when 16#0B8D# => romdata <= X"F068A6CA";
    when 16#0B8E# => romdata <= X"1442AF77";
    when 16#0B8F# => romdata <= X"C83B7D86";
    when 16#0B90# => romdata <= X"49DC281B";
    when 16#0B91# => romdata <= X"F438F957";
    when 16#0B92# => romdata <= X"6F7A719A";
    when 16#0B93# => romdata <= X"902A860B";
    when 16#0B94# => romdata <= X"9ECE9AE9";
    when 16#0B95# => romdata <= X"C14B9885";
    when 16#0B96# => romdata <= X"9B282010";
    when 16#0B97# => romdata <= X"A5DC90DC";
    when 16#0B98# => romdata <= X"E612AFEF";
    when 16#0B99# => romdata <= X"D44E0E9E";
    when 16#0B9A# => romdata <= X"7666A461";
    when 16#0B9B# => romdata <= X"AE50C265";
    when 16#0B9C# => romdata <= X"6BC03664";
    when 16#0B9D# => romdata <= X"8B826CA9";
    when 16#0B9E# => romdata <= X"C3C7C53B";
    when 16#0B9F# => romdata <= X"30976335";
    when 16#0BA0# => romdata <= X"B097C193";
    when 16#0BA1# => romdata <= X"90716A41";
    when 16#0BA2# => romdata <= X"FD437A20";
    when 16#0BA3# => romdata <= X"98BCFA2B";
    when 16#0BA4# => romdata <= X"2975F1EA";
    when 16#0BA5# => romdata <= X"E5BDBB81";
    when 16#0BA6# => romdata <= X"92024C20";
    when 16#0BA7# => romdata <= X"136D2542";
    when 16#0BA8# => romdata <= X"FD89FB8F";
    when 16#0BA9# => romdata <= X"2F94C08F";
    when 16#0BAA# => romdata <= X"76510927";
    when 16#0BAB# => romdata <= X"9BC4E511";
    when 16#0BAC# => romdata <= X"78749623";
    when 16#0BAD# => romdata <= X"3F15F52D";
    when 16#0BAE# => romdata <= X"7C3BC3E9";
    when 16#0BAF# => romdata <= X"8A6DC39A";
    when 16#0BB0# => romdata <= X"FA1818B9";
    when 16#0BB1# => romdata <= X"533EDE72";
    when 16#0BB2# => romdata <= X"FDAF021E";
    when 16#0BB3# => romdata <= X"2C9B7D6C";
    when 16#0BB4# => romdata <= X"74E49B84";
    when 16#0BB5# => romdata <= X"9F372B1A";
    when 16#0BB6# => romdata <= X"131F4C53";
    when 16#0BB7# => romdata <= X"2DBE3B63";
    when 16#0BB8# => romdata <= X"635E0E13";
    when 16#0BB9# => romdata <= X"34C87DDB";
    when 16#0BBA# => romdata <= X"6F3D7388";
    when 16#0BBB# => romdata <= X"3D2B43E8";
    when 16#0BBC# => romdata <= X"7CF19E40";
    when 16#0BBD# => romdata <= X"D6B404E5";
    when 16#0BBE# => romdata <= X"81E807E6";
    when 16#0BBF# => romdata <= X"EC1A94F5";
    when 16#0BC0# => romdata <= X"261C7F7E";
    when 16#0BC1# => romdata <= X"FD4CF043";
    when 16#0BC2# => romdata <= X"C90A1A7E";
    when 16#0BC3# => romdata <= X"97465022";
    when 16#0BC4# => romdata <= X"ABAA1DC2";
    when 16#0BC5# => romdata <= X"1588FD28";
    when 16#0BC6# => romdata <= X"5E7158FD";
    when 16#0BC7# => romdata <= X"9B67EC5F";
    when 16#0BC8# => romdata <= X"E7C9E840";
    when 16#0BC9# => romdata <= X"29E961E0";
    when 16#0BCA# => romdata <= X"45EB5227";
    when 16#0BCB# => romdata <= X"E4726154";
    when 16#0BCC# => romdata <= X"F4F057FA";
    when 16#0BCD# => romdata <= X"337BB20D";
    when 16#0BCE# => romdata <= X"DA25D116";
    when 16#0BCF# => romdata <= X"32A7995B";
    when 16#0BD0# => romdata <= X"81076408";
    when 16#0BD1# => romdata <= X"4EBDE01A";
    when 16#0BD2# => romdata <= X"F07372EA";
    when 16#0BD3# => romdata <= X"82FBAFE0";
    when 16#0BD4# => romdata <= X"434401FC";
    when 16#0BD5# => romdata <= X"FE05CE8F";
    when 16#0BD6# => romdata <= X"E3C20C01";
    when 16#0BD7# => romdata <= X"ACF4E9B8";
    when 16#0BD8# => romdata <= X"EAF4D50C";
    when 16#0BD9# => romdata <= X"73D5C42A";
    when 16#0BDA# => romdata <= X"95526CDC";
    when 16#0BDB# => romdata <= X"8313DBCA";
    when 16#0BDC# => romdata <= X"6ECEACB4";
    when 16#0BDD# => romdata <= X"57D96735";
    when 16#0BDE# => romdata <= X"65A1CC0A";
    when 16#0BDF# => romdata <= X"AE23FD62";
    when 16#0BE0# => romdata <= X"61A8943E";
    when 16#0BE1# => romdata <= X"8FB84CCE";
    when 16#0BE2# => romdata <= X"C676601A";
    when 16#0BE3# => romdata <= X"4B302A9C";
    when 16#0BE4# => romdata <= X"ACDEC899";
    when 16#0BE5# => romdata <= X"8EDC847A";
    when 16#0BE6# => romdata <= X"53B3CB0E";
    when 16#0BE7# => romdata <= X"12C8B4A7";
    when 16#0BE8# => romdata <= X"897D5680";
    when 16#0BE9# => romdata <= X"CB14A3D1";
    when 16#0BEA# => romdata <= X"1BDBF482";
    when 16#0BEB# => romdata <= X"6C3938EB";
    when 16#0BEC# => romdata <= X"EEFA0075";
    when 16#0BED# => romdata <= X"B6494CC7";
    when 16#0BEE# => romdata <= X"14D3C0DD";
    when 16#0BEF# => romdata <= X"A2F5F783";
    when 16#0BF0# => romdata <= X"CF23AD2D";
    when 16#0BF1# => romdata <= X"2545C899";
    when 16#0BF2# => romdata <= X"867C1115";
    when 16#0BF3# => romdata <= X"BF4A4F55";
    when 16#0BF4# => romdata <= X"9F63E680";
    when 16#0BF5# => romdata <= X"98955550";
    when 16#0BF6# => romdata <= X"BFA1EF77";
    when 16#0BF7# => romdata <= X"71598EF8";
    when 16#0BF8# => romdata <= X"6A08C0C6";
    when 16#0BF9# => romdata <= X"34B29167";
    when 16#0BFA# => romdata <= X"4BB77615";
    when 16#0BFB# => romdata <= X"121BF083";
    when 16#0BFC# => romdata <= X"8DA96D6E";
    when 16#0BFD# => romdata <= X"7C53BFE6";
    when 16#0BFE# => romdata <= X"A58A382F";
    when 16#0BFF# => romdata <= X"D9721CC0";
    when 16#0C00# => romdata <= X"BF8903A3";
    when 16#0C01# => romdata <= X"918B3FDC";
    when 16#0C02# => romdata <= X"06CAB4EF";
    when 16#0C03# => romdata <= X"675F7BE3";
    when 16#0C04# => romdata <= X"962CD7E3";
    when 16#0C05# => romdata <= X"C6ED6433";
    when 16#0C06# => romdata <= X"86EE533C";
    when 16#0C07# => romdata <= X"3B24A3D9";
    when 16#0C08# => romdata <= X"4D2EA2CF";
    when 16#0C09# => romdata <= X"B83F0A34";
    when 16#0C0A# => romdata <= X"6FF2875D";
    when 16#0C0B# => romdata <= X"B07BA647";
    when 16#0C0C# => romdata <= X"492D47A8";
    when 16#0C0D# => romdata <= X"07E7FD97";
    when 16#0C0E# => romdata <= X"17CF12BC";
    when 16#0C0F# => romdata <= X"97B3C1BE";
    when 16#0C10# => romdata <= X"1361E598";
    when 16#0C11# => romdata <= X"850B39D5";
    when 16#0C12# => romdata <= X"0CF7BE70";
    when 16#0C13# => romdata <= X"0507863B";
    when 16#0C14# => romdata <= X"C4BBF266";
    when 16#0C15# => romdata <= X"20FAC11D";
    when 16#0C16# => romdata <= X"97128049";
    when 16#0C17# => romdata <= X"BD96C5E0";
    when 16#0C18# => romdata <= X"9DC8FF3F";
    when 16#0C19# => romdata <= X"62655D66";
    when 16#0C1A# => romdata <= X"0FE66D31";
    when 16#0C1B# => romdata <= X"AB0B0F6D";
    when 16#0C1C# => romdata <= X"4F8420E3";
    when 16#0C1D# => romdata <= X"D2E633C5";
    when 16#0C1E# => romdata <= X"71D7FE2A";
    when 16#0C1F# => romdata <= X"F1CB4E3B";
    when 16#0C20# => romdata <= X"EE95E092";
    when 16#0C21# => romdata <= X"B00EFD27";
    when 16#0C22# => romdata <= X"96A3DEF3";
    when 16#0C23# => romdata <= X"76F75B7E";
    when 16#0C24# => romdata <= X"FCBB1413";
    when 16#0C25# => romdata <= X"37D81AE5";
    when 16#0C26# => romdata <= X"2939D879";
    when 16#0C27# => romdata <= X"56C41B1E";
    when 16#0C28# => romdata <= X"42C1CCA4";
    when 16#0C29# => romdata <= X"317D31AB";
    when 16#0C2A# => romdata <= X"4F53DC95";
    when 16#0C2B# => romdata <= X"02A3DC77";
    when 16#0C2C# => romdata <= X"4E05E1ED";
    when 16#0C2D# => romdata <= X"5008CD93";
    when 16#0C2E# => romdata <= X"1DDDB98D";
    when 16#0C2F# => romdata <= X"FA69960A";
    when 16#0C30# => romdata <= X"6ACD45B6";
    when 16#0C31# => romdata <= X"0895C4FB";
    when 16#0C32# => romdata <= X"A2BDAE8B";
    when 16#0C33# => romdata <= X"C7DB8C82";
    when 16#0C34# => romdata <= X"1697558B";
    when 16#0C35# => romdata <= X"1E0A3111";
    when 16#0C36# => romdata <= X"F1567384";
    when 16#0C37# => romdata <= X"09FD180C";
    when 16#0C38# => romdata <= X"5A4A33B2";
    when 16#0C39# => romdata <= X"4C5EE499";
    when 16#0C3A# => romdata <= X"1B84133C";
    when 16#0C3B# => romdata <= X"E9AC0897";
    when 16#0C3C# => romdata <= X"24D62DA9";
    when 16#0C3D# => romdata <= X"D9827A2A";
    when 16#0C3E# => romdata <= X"04FC1036";
    when 16#0C3F# => romdata <= X"52F216A0";
    when 16#0C40# => romdata <= X"895E78A9";
    when 16#0C41# => romdata <= X"60862708";
    when 16#0C42# => romdata <= X"14C2699F";
    when 16#0C43# => romdata <= X"475CEFD6";
    when 16#0C44# => romdata <= X"359428D8";
    when 16#0C45# => romdata <= X"C505BBE8";
    when 16#0C46# => romdata <= X"C1A96D27";
    when 16#0C47# => romdata <= X"93802219";
    when 16#0C48# => romdata <= X"144CA6B3";
    when 16#0C49# => romdata <= X"EDB45592";
    when 16#0C4A# => romdata <= X"9B39A3E9";
    when 16#0C4B# => romdata <= X"F3AB74D6";
    when 16#0C4C# => romdata <= X"85608CE3";
    when 16#0C4D# => romdata <= X"F301FE38";
    when 16#0C4E# => romdata <= X"202ADFEF";
    when 16#0C4F# => romdata <= X"529CCFF4";
    when 16#0C50# => romdata <= X"6AF36DC2";
    when 16#0C51# => romdata <= X"4956A7CD";
    when 16#0C52# => romdata <= X"07CEBA55";
    when 16#0C53# => romdata <= X"AA4C89F7";
    when 16#0C54# => romdata <= X"913A8A4B";
    when 16#0C55# => romdata <= X"844FD8F1";
    when 16#0C56# => romdata <= X"52C8A823";
    when 16#0C57# => romdata <= X"CB9888E3";
    when 16#0C58# => romdata <= X"BFEA97D7";
    when 16#0C59# => romdata <= X"E4AAFA07";
    when 16#0C5A# => romdata <= X"125DA4F5";
    when 16#0C5B# => romdata <= X"1D974A5D";
    when 16#0C5C# => romdata <= X"AFF0045B";
    when 16#0C5D# => romdata <= X"CE5B8681";
    when 16#0C5E# => romdata <= X"77A91BD9";
    when 16#0C5F# => romdata <= X"32963451";
    when 16#0C60# => romdata <= X"EE2673A8";
    when 16#0C61# => romdata <= X"5AA8B7D4";
    when 16#0C62# => romdata <= X"93BDF25B";
    when 16#0C63# => romdata <= X"CC2F64AE";
    when 16#0C64# => romdata <= X"C3150D8C";
    when 16#0C65# => romdata <= X"40C835AB";
    when 16#0C66# => romdata <= X"4F5D0B7F";
    when 16#0C67# => romdata <= X"259DF099";
    when 16#0C68# => romdata <= X"BD6FA9F5";
    when 16#0C69# => romdata <= X"CB198B61";
    when 16#0C6A# => romdata <= X"018B1448";
    when 16#0C6B# => romdata <= X"035CCD34";
    when 16#0C6C# => romdata <= X"E7E7A213";
    when 16#0C6D# => romdata <= X"8F437490";
    when 16#0C6E# => romdata <= X"026050BB";
    when 16#0C6F# => romdata <= X"E3CE2D4C";
    when 16#0C70# => romdata <= X"F4F4F095";
    when 16#0C71# => romdata <= X"CB97548E";
    when 16#0C72# => romdata <= X"5731A338";
    when 16#0C73# => romdata <= X"CB390351";
    when 16#0C74# => romdata <= X"9D6B13A0";
    when 16#0C75# => romdata <= X"29727F04";
    when 16#0C76# => romdata <= X"7A7D0090";
    when 16#0C77# => romdata <= X"4A556C88";
    when 16#0C78# => romdata <= X"37454103";
    when 16#0C79# => romdata <= X"60FC878F";
    when 16#0C7A# => romdata <= X"77707A71";
    when 16#0C7B# => romdata <= X"6D549ACD";
    when 16#0C7C# => romdata <= X"6A70A18F";
    when 16#0C7D# => romdata <= X"9EE0AA8A";
    when 16#0C7E# => romdata <= X"6EE20806";
    when 16#0C7F# => romdata <= X"08E10AC0";
    when 16#0C80# => romdata <= X"F58CDE0E";
    when 16#0C81# => romdata <= X"FE2356F4";
    when 16#0C82# => romdata <= X"29B0F2F9";
    when 16#0C83# => romdata <= X"A7869A41";
    when 16#0C84# => romdata <= X"42A61731";
    when 16#0C85# => romdata <= X"88DD75B5";
    when 16#0C86# => romdata <= X"70F1D1EC";
    when 16#0C87# => romdata <= X"D282E4AF";
    when 16#0C88# => romdata <= X"BAD11370";
    when 16#0C89# => romdata <= X"C5B4CCF3";
    when 16#0C8A# => romdata <= X"C98535D2";
    when 16#0C8B# => romdata <= X"7D73C011";
    when 16#0C8C# => romdata <= X"1F11A847";
    when 16#0C8D# => romdata <= X"11F73244";
    when 16#0C8E# => romdata <= X"1EAECAB6";
    when 16#0C8F# => romdata <= X"84F2F0D7";
    when 16#0C90# => romdata <= X"FD4FC407";
    when 16#0C91# => romdata <= X"07495749";
    when 16#0C92# => romdata <= X"22A906E8";
    when 16#0C93# => romdata <= X"4B3350CD";
    when 16#0C94# => romdata <= X"E5957DC3";
    when 16#0C95# => romdata <= X"88FDA23B";
    when 16#0C96# => romdata <= X"F45F0595";
    when 16#0C97# => romdata <= X"1A393DA2";
    when 16#0C98# => romdata <= X"53EAF691";
    when 16#0C99# => romdata <= X"940897B5";
    when 16#0C9A# => romdata <= X"7ACE655E";
    when 16#0C9B# => romdata <= X"9630F098";
    when 16#0C9C# => romdata <= X"56E76958";
    when 16#0C9D# => romdata <= X"D6BF7B83";
    when 16#0C9E# => romdata <= X"0E0CB818";
    when 16#0C9F# => romdata <= X"2AE226F3";
    when 16#0CA0# => romdata <= X"9D48036C";
    when 16#0CA1# => romdata <= X"867BEFA7";
    when 16#0CA2# => romdata <= X"E7ADBAD1";
    when 16#0CA3# => romdata <= X"7C1AB452";
    when 16#0CA4# => romdata <= X"97C757DA";
    when 16#0CA5# => romdata <= X"4AFFBAE6";
    when 16#0CA6# => romdata <= X"77B05677";
    when 16#0CA7# => romdata <= X"D60DE1D9";
    when 16#0CA8# => romdata <= X"75A4F3D7";
    when 16#0CA9# => romdata <= X"EB3461B4";
    when 16#0CAA# => romdata <= X"24B67B61";
    when 16#0CAB# => romdata <= X"025AAC25";
    when 16#0CAC# => romdata <= X"7A69FF72";
    when 16#0CAD# => romdata <= X"0CB9DAC0";
    when 16#0CAE# => romdata <= X"07C50C69";
    when 16#0CAF# => romdata <= X"A7ACDBBC";
    when 16#0CB0# => romdata <= X"E210BAD4";
    when 16#0CB1# => romdata <= X"DC2E629A";
    when 16#0CB2# => romdata <= X"039D98E7";
    when 16#0CB3# => romdata <= X"EA037A5C";
    when 16#0CB4# => romdata <= X"344B5CAE";
    when 16#0CB5# => romdata <= X"DCDA035F";
    when 16#0CB6# => romdata <= X"28677A41";
    when 16#0CB7# => romdata <= X"D55A0E3E";
    when 16#0CB8# => romdata <= X"6E480CCB";
    when 16#0CB9# => romdata <= X"12B8F170";
    when 16#0CBA# => romdata <= X"62A983F4";
    when 16#0CBB# => romdata <= X"E651B4F7";
    when 16#0CBC# => romdata <= X"CB217FD0";
    when 16#0CBD# => romdata <= X"6BE46747";
    when 16#0CBE# => romdata <= X"CD5418C0";
    when 16#0CBF# => romdata <= X"C8191646";
    when 16#0CC0# => romdata <= X"5A4F5660";
    when 16#0CC1# => romdata <= X"152B3E47";
    when 16#0CC2# => romdata <= X"81DA8040";
    when 16#0CC3# => romdata <= X"D4246F9B";
    when 16#0CC4# => romdata <= X"C47366BF";
    when 16#0CC5# => romdata <= X"663CF9DA";
    when 16#0CC6# => romdata <= X"3BB247D9";
    when 16#0CC7# => romdata <= X"238873CC";
    when 16#0CC8# => romdata <= X"DC6FC62D";
    when 16#0CC9# => romdata <= X"1D8F669E";
    when 16#0CCA# => romdata <= X"FBA42527";
    when 16#0CCB# => romdata <= X"112FF407";
    when 16#0CCC# => romdata <= X"2262F7E6";
    when 16#0CCD# => romdata <= X"5AEAC328";
    when 16#0CCE# => romdata <= X"871DDF47";
    when 16#0CCF# => romdata <= X"588A0A0D";
    when 16#0CD0# => romdata <= X"D13A4139";
    when 16#0CD1# => romdata <= X"F4145822";
    when 16#0CD2# => romdata <= X"A5917F62";
    when 16#0CD3# => romdata <= X"4B881BFC";
    when 16#0CD4# => romdata <= X"354F37B6";
    when 16#0CD5# => romdata <= X"D59C5668";
    when 16#0CD6# => romdata <= X"23F629A2";
    when 16#0CD7# => romdata <= X"1C973324";
    when 16#0CD8# => romdata <= X"F7167BC3";
    when 16#0CD9# => romdata <= X"9FBD2C12";
    when 16#0CDA# => romdata <= X"1D2A8493";
    when 16#0CDB# => romdata <= X"08D13DA1";
    when 16#0CDC# => romdata <= X"A28948EB";
    when 16#0CDD# => romdata <= X"59F7DE97";
    when 16#0CDE# => romdata <= X"E364223E";
    when 16#0CDF# => romdata <= X"17A30119";
    when 16#0CE0# => romdata <= X"BBC7F43E";
    when 16#0CE1# => romdata <= X"21E7DC30";
    when 16#0CE2# => romdata <= X"93F75050";
    when 16#0CE3# => romdata <= X"55ADAB46";
    when 16#0CE4# => romdata <= X"54194A77";
    when 16#0CE5# => romdata <= X"C1CCB618";
    when 16#0CE6# => romdata <= X"98840125";
    when 16#0CE7# => romdata <= X"455A275A";
    when 16#0CE8# => romdata <= X"8F071273";
    when 16#0CE9# => romdata <= X"D8C13934";
    when 16#0CEA# => romdata <= X"915D379C";
    when 16#0CEB# => romdata <= X"C603657D";
    when 16#0CEC# => romdata <= X"99CE4075";
    when 16#0CED# => romdata <= X"C1F1DCAB";
    when 16#0CEE# => romdata <= X"60B6BD62";
    when 16#0CEF# => romdata <= X"ABA1A10B";
    when 16#0CF0# => romdata <= X"5402A597";
    when 16#0CF1# => romdata <= X"06798002";
    when 16#0CF2# => romdata <= X"EF30ADED";
    when 16#0CF3# => romdata <= X"2F354E38";
    when 16#0CF4# => romdata <= X"CE0B5790";
    when 16#0CF5# => romdata <= X"0FDAD31E";
    when 16#0CF6# => romdata <= X"7F684E53";
    when 16#0CF7# => romdata <= X"D097B431";
    when 16#0CF8# => romdata <= X"3DB552EA";
    when 16#0CF9# => romdata <= X"66F6D337";
    when 16#0CFA# => romdata <= X"F2959447";
    when 16#0CFB# => romdata <= X"0D3DC0BC";
    when 16#0CFC# => romdata <= X"6CD36183";
    when 16#0CFD# => romdata <= X"1251004D";
    when 16#0CFE# => romdata <= X"D3C5357B";
    when 16#0CFF# => romdata <= X"C0BECFE0";
    when 16#0D00# => romdata <= X"D9086F7C";
    when 16#0D01# => romdata <= X"272AA317";
    when 16#0D02# => romdata <= X"C64C00AF";
    when 16#0D03# => romdata <= X"43C924DB";
    when 16#0D04# => romdata <= X"5DAC97F8";
    when 16#0D05# => romdata <= X"EE3ED229";
    when 16#0D06# => romdata <= X"6252FC47";
    when 16#0D07# => romdata <= X"56FCE692";
    when 16#0D08# => romdata <= X"8BB009D4";
    when 16#0D09# => romdata <= X"488B9BAB";
    when 16#0D0A# => romdata <= X"757411BB";
    when 16#0D0B# => romdata <= X"A52BA6F6";
    when 16#0D0C# => romdata <= X"1AF1181C";
    when 16#0D0D# => romdata <= X"C7BBA942";
    when 16#0D0E# => romdata <= X"57593FA1";
    when 16#0D0F# => romdata <= X"BD26D52A";
    when 16#0D10# => romdata <= X"D5014C3F";
    when 16#0D11# => romdata <= X"1A1832FC";
    when 16#0D12# => romdata <= X"4F7445C8";
    when 16#0D13# => romdata <= X"BBB77C8F";
    when 16#0D14# => romdata <= X"D31C88F0";
    when 16#0D15# => romdata <= X"C5D4736D";
    when 16#0D16# => romdata <= X"49DCDFBE";
    when 16#0D17# => romdata <= X"EF2B8301";
    when 16#0D18# => romdata <= X"E3118579";
    when 16#0D19# => romdata <= X"3BFF87CF";
    when 16#0D1A# => romdata <= X"D9E6F7E0";
    when 16#0D1B# => romdata <= X"84D343AB";
    when 16#0D1C# => romdata <= X"98BA3518";
    when 16#0D1D# => romdata <= X"A87A5F91";
    when 16#0D1E# => romdata <= X"5BC0D76B";
    when 16#0D1F# => romdata <= X"01AF7DC1";
    when 16#0D20# => romdata <= X"CE45F1C5";
    when 16#0D21# => romdata <= X"280BD39D";
    when 16#0D22# => romdata <= X"3E3D94D0";
    when 16#0D23# => romdata <= X"A0286F8B";
    when 16#0D24# => romdata <= X"D9FA9428";
    when 16#0D25# => romdata <= X"49664E08";
    when 16#0D26# => romdata <= X"F2BE0B93";
    when 16#0D27# => romdata <= X"C6E3B890";
    when 16#0D28# => romdata <= X"61193FAD";
    when 16#0D29# => romdata <= X"A0FA9485";
    when 16#0D2A# => romdata <= X"F62CA87F";
    when 16#0D2B# => romdata <= X"3E68E204";
    when 16#0D2C# => romdata <= X"186EF118";
    when 16#0D2D# => romdata <= X"7642D651";
    when 16#0D2E# => romdata <= X"162E4D8E";
    when 16#0D2F# => romdata <= X"7DA049F4";
    when 16#0D30# => romdata <= X"62362D8C";
    when 16#0D31# => romdata <= X"94539CAA";
    when 16#0D32# => romdata <= X"D09AE476";
    when 16#0D33# => romdata <= X"8C96ED6C";
    when 16#0D34# => romdata <= X"2CAB8025";
    when 16#0D35# => romdata <= X"EBB6901C";
    when 16#0D36# => romdata <= X"BB26865E";
    when 16#0D37# => romdata <= X"1F19FA1B";
    when 16#0D38# => romdata <= X"193D47EC";
    when 16#0D39# => romdata <= X"E390B881";
    when 16#0D3A# => romdata <= X"23357895";
    when 16#0D3B# => romdata <= X"0175C85B";
    when 16#0D3C# => romdata <= X"928582D5";
    when 16#0D3D# => romdata <= X"B439EEF2";
    when 16#0D3E# => romdata <= X"F56A8C7E";
    when 16#0D3F# => romdata <= X"A09278E4";
    when 16#0D40# => romdata <= X"77410512";
    when 16#0D41# => romdata <= X"23AC1824";
    when 16#0D42# => romdata <= X"56C4FA04";
    when 16#0D43# => romdata <= X"D025BDB3";
    when 16#0D44# => romdata <= X"3FA10C48";
    when 16#0D45# => romdata <= X"C70EC91B";
    when 16#0D46# => romdata <= X"C709E3CB";
    when 16#0D47# => romdata <= X"0FA3E01D";
    when 16#0D48# => romdata <= X"CE5FE5EC";
    when 16#0D49# => romdata <= X"B9018130";
    when 16#0D4A# => romdata <= X"A8DE5D05";
    when 16#0D4B# => romdata <= X"83EDD68E";
    when 16#0D4C# => romdata <= X"A2EF227A";
    when 16#0D4D# => romdata <= X"612748B2";
    when 16#0D4E# => romdata <= X"F785A30A";
    when 16#0D4F# => romdata <= X"01014BD4";
    when 16#0D50# => romdata <= X"79DEC625";
    when 16#0D51# => romdata <= X"6C8AD884";
    when 16#0D52# => romdata <= X"70F79DE0";
    when 16#0D53# => romdata <= X"E1432CAE";
    when 16#0D54# => romdata <= X"448DD704";
    when 16#0D55# => romdata <= X"9E5B7D4D";
    when 16#0D56# => romdata <= X"F3C978F6";
    when 16#0D57# => romdata <= X"5E708CA3";
    when 16#0D58# => romdata <= X"759AAB9D";
    when 16#0D59# => romdata <= X"329C11FA";
    when 16#0D5A# => romdata <= X"D71204E1";
    when 16#0D5B# => romdata <= X"E92322E3";
    when 16#0D5C# => romdata <= X"EA1BBDD9";
    when 16#0D5D# => romdata <= X"D034E2A2";
    when 16#0D5E# => romdata <= X"3ACAFA21";
    when 16#0D5F# => romdata <= X"CF490AA5";
    when 16#0D60# => romdata <= X"E2E41919";
    when 16#0D61# => romdata <= X"7DBE9906";
    when 16#0D62# => romdata <= X"67BCF277";
    when 16#0D63# => romdata <= X"ED61B264";
    when 16#0D64# => romdata <= X"632F6943";
    when 16#0D65# => romdata <= X"92EF52F0";
    when 16#0D66# => romdata <= X"A27C38E4";
    when 16#0D67# => romdata <= X"78257AEC";
    when 16#0D68# => romdata <= X"8D254293";
    when 16#0D69# => romdata <= X"8BF0713E";
    when 16#0D6A# => romdata <= X"BE60779C";
    when 16#0D6B# => romdata <= X"95A0EEC8";
    when 16#0D6C# => romdata <= X"F32A5202";
    when 16#0D6D# => romdata <= X"A849CEE8";
    when 16#0D6E# => romdata <= X"CE0F9970";
    when 16#0D6F# => romdata <= X"2F595AEA";
    when 16#0D70# => romdata <= X"839531D4";
    when 16#0D71# => romdata <= X"CFB5F5A6";
    when 16#0D72# => romdata <= X"166B06EB";
    when 16#0D73# => romdata <= X"64387552";
    when 16#0D74# => romdata <= X"A1F9BC6B";
    when 16#0D75# => romdata <= X"B97B9B99";
    when 16#0D76# => romdata <= X"D19C3D2E";
    when 16#0D77# => romdata <= X"1E8E9B30";
    when 16#0D78# => romdata <= X"5D525E74";
    when 16#0D79# => romdata <= X"13496E40";
    when 16#0D7A# => romdata <= X"FF50CF77";
    when 16#0D7B# => romdata <= X"D4D4E2D4";
    when 16#0D7C# => romdata <= X"1B1D5929";
    when 16#0D7D# => romdata <= X"848FB2F1";
    when 16#0D7E# => romdata <= X"FDDA5A39";
    when 16#0D7F# => romdata <= X"DEA05460";
    when 16#0D80# => romdata <= X"AE4E3B30";
    when 16#0D81# => romdata <= X"560A50DA";
    when 16#0D82# => romdata <= X"55AB3E59";
    when 16#0D83# => romdata <= X"FFF51284";
    when 16#0D84# => romdata <= X"4A2700D2";
    when 16#0D85# => romdata <= X"D763D85D";
    when 16#0D86# => romdata <= X"5C3FD8CF";
    when 16#0D87# => romdata <= X"EFACD4D0";
    when 16#0D88# => romdata <= X"23BD926D";
    when 16#0D89# => romdata <= X"3EF2E55E";
    when 16#0D8A# => romdata <= X"B1B3831F";
    when 16#0D8B# => romdata <= X"2276EB07";
    when 16#0D8C# => romdata <= X"E5C07B44";
    when 16#0D8D# => romdata <= X"FD7D7933";
    when 16#0D8E# => romdata <= X"3699BED0";
    when 16#0D8F# => romdata <= X"804B6789";
    when 16#0D90# => romdata <= X"15FE0F09";
    when 16#0D91# => romdata <= X"2DA9A62F";
    when 16#0D92# => romdata <= X"69CB020D";
    when 16#0D93# => romdata <= X"A21932F9";
    when 16#0D94# => romdata <= X"FDF9AF33";
    when 16#0D95# => romdata <= X"2E1B400C";
    when 16#0D96# => romdata <= X"6B7E7880";
    when 16#0D97# => romdata <= X"508E840D";
    when 16#0D98# => romdata <= X"62FBA07E";
    when 16#0D99# => romdata <= X"827A23A2";
    when 16#0D9A# => romdata <= X"575AE68E";
    when 16#0D9B# => romdata <= X"15AC444A";
    when 16#0D9C# => romdata <= X"1CE35DF3";
    when 16#0D9D# => romdata <= X"C3F7CA49";
    when 16#0D9E# => romdata <= X"DEF2966D";
    when 16#0D9F# => romdata <= X"F3BA89C8";
    when 16#0DA0# => romdata <= X"E90ED5E2";
    when 16#0DA1# => romdata <= X"421A6407";
    when 16#0DA2# => romdata <= X"F2EC51A3";
    when 16#0DA3# => romdata <= X"E92A3608";
    when 16#0DA4# => romdata <= X"FCBD6AD9";
    when 16#0DA5# => romdata <= X"FF9E5C78";
    when 16#0DA6# => romdata <= X"17E79A0C";
    when 16#0DA7# => romdata <= X"09FE9014";
    when 16#0DA8# => romdata <= X"F7AC2914";
    when 16#0DA9# => romdata <= X"48263E43";
    when 16#0DAA# => romdata <= X"46CBC4BA";
    when 16#0DAB# => romdata <= X"A6EABFB5";
    when 16#0DAC# => romdata <= X"9B4526B6";
    when 16#0DAD# => romdata <= X"54070084";
    when 16#0DAE# => romdata <= X"F52B864F";
    when 16#0DAF# => romdata <= X"9769181D";
    when 16#0DB0# => romdata <= X"C6EA91B5";
    when 16#0DB1# => romdata <= X"76956397";
    when 16#0DB2# => romdata <= X"CE55CCDD";
    when 16#0DB3# => romdata <= X"BE41F94E";
    when 16#0DB4# => romdata <= X"5DC366E7";
    when 16#0DB5# => romdata <= X"75C86ADB";
    when 16#0DB6# => romdata <= X"1C807B66";
    when 16#0DB7# => romdata <= X"D08696A2";
    when 16#0DB8# => romdata <= X"BEE45B90";
    when 16#0DB9# => romdata <= X"E8736469";
    when 16#0DBA# => romdata <= X"A371F059";
    when 16#0DBB# => romdata <= X"29D9D9FD";
    when 16#0DBC# => romdata <= X"34980DE0";
    when 16#0DBD# => romdata <= X"8E00BDE2";
    when 16#0DBE# => romdata <= X"CD0EAB6A";
    when 16#0DBF# => romdata <= X"F2165D76";
    when 16#0DC0# => romdata <= X"519F8F2D";
    when 16#0DC1# => romdata <= X"894AC707";
    when 16#0DC2# => romdata <= X"40D2372B";
    when 16#0DC3# => romdata <= X"37407BDA";
    when 16#0DC4# => romdata <= X"4D943EDF";
    when 16#0DC5# => romdata <= X"1CBD35CC";
    when 16#0DC6# => romdata <= X"E4D81340";
    when 16#0DC7# => romdata <= X"CC97751C";
    when 16#0DC8# => romdata <= X"568731C0";
    when 16#0DC9# => romdata <= X"09DF6557";
    when 16#0DCA# => romdata <= X"1F28B7F5";
    when 16#0DCB# => romdata <= X"8106AE67";
    when 16#0DCC# => romdata <= X"279E83C3";
    when 16#0DCD# => romdata <= X"A0C130DE";
    when 16#0DCE# => romdata <= X"0C5B6C99";
    when 16#0DCF# => romdata <= X"11709954";
    when 16#0DD0# => romdata <= X"8661D290";
    when 16#0DD1# => romdata <= X"C4CAF3BC";
    when 16#0DD2# => romdata <= X"60EF719E";
    when 16#0DD3# => romdata <= X"2F7B210F";
    when 16#0DD4# => romdata <= X"CD4381C3";
    when 16#0DD5# => romdata <= X"3904AFDF";
    when 16#0DD6# => romdata <= X"96DC3A65";
    when 16#0DD7# => romdata <= X"57B42B6E";
    when 16#0DD8# => romdata <= X"E895B4D6";
    when 16#0DD9# => romdata <= X"04F5F898";
    when 16#0DDA# => romdata <= X"5F454C51";
    when 16#0DDB# => romdata <= X"E32B2C87";
    when 16#0DDC# => romdata <= X"4E90926C";
    when 16#0DDD# => romdata <= X"BC58D044";
    when 16#0DDE# => romdata <= X"D483D6D2";
    when 16#0DDF# => romdata <= X"A7C26C7A";
    when 16#0DE0# => romdata <= X"C4D19053";
    when 16#0DE1# => romdata <= X"1F79993D";
    when 16#0DE2# => romdata <= X"07B2E830";
    when 16#0DE3# => romdata <= X"FEB99BFD";
    when 16#0DE4# => romdata <= X"B00AE8C0";
    when 16#0DE5# => romdata <= X"08DB1B76";
    when 16#0DE6# => romdata <= X"2F3F4A81";
    when 16#0DE7# => romdata <= X"D41295FD";
    when 16#0DE8# => romdata <= X"DA37F305";
    when 16#0DE9# => romdata <= X"6B1110D4";
    when 16#0DEA# => romdata <= X"F0CF385F";
    when 16#0DEB# => romdata <= X"9FCC7E14";
    when 16#0DEC# => romdata <= X"C34F6752";
    when 16#0DED# => romdata <= X"A2FB17F5";
    when 16#0DEE# => romdata <= X"CD3FC4AF";
    when 16#0DEF# => romdata <= X"0D51E4A0";
    when 16#0DF0# => romdata <= X"AF7D28DB";
    when 16#0DF1# => romdata <= X"0D4D6511";
    when 16#0DF2# => romdata <= X"56189209";
    when 16#0DF3# => romdata <= X"480054F8";
    when 16#0DF4# => romdata <= X"287266B1";
    when 16#0DF5# => romdata <= X"CB26C9E8";
    when 16#0DF6# => romdata <= X"CACAA0BE";
    when 16#0DF7# => romdata <= X"5A69C696";
    when 16#0DF8# => romdata <= X"300025D1";
    when 16#0DF9# => romdata <= X"60F9DA29";
    when 16#0DFA# => romdata <= X"F9EC7983";
    when 16#0DFB# => romdata <= X"8941459B";
    when 16#0DFC# => romdata <= X"7B8164AA";
    when 16#0DFD# => romdata <= X"D95577A0";
    when 16#0DFE# => romdata <= X"C532EC2E";
    when 16#0DFF# => romdata <= X"DB352500";
    when 16#0E00# => romdata <= X"9CF0CC00";
    when 16#0E01# => romdata <= X"B5788DD7";
    when 16#0E02# => romdata <= X"43A5F33D";
    when 16#0E03# => romdata <= X"87E8FA57";
    when 16#0E04# => romdata <= X"33B72EDB";
    when 16#0E05# => romdata <= X"CD61AA4B";
    when 16#0E06# => romdata <= X"8D0B8121";
    when 16#0E07# => romdata <= X"3DB52E7E";
    when 16#0E08# => romdata <= X"F17AE909";
    when 16#0E09# => romdata <= X"34F5EC07";
    when 16#0E0A# => romdata <= X"11ADD19E";
    when 16#0E0B# => romdata <= X"881CC330";
    when 16#0E0C# => romdata <= X"F696179C";
    when 16#0E0D# => romdata <= X"1BA464FF";
    when 16#0E0E# => romdata <= X"E6D7B04E";
    when 16#0E0F# => romdata <= X"EC383A41";
    when 16#0E10# => romdata <= X"06BE5892";
    when 16#0E11# => romdata <= X"C5DD1BD7";
    when 16#0E12# => romdata <= X"19AB3739";
    when 16#0E13# => romdata <= X"A909A384";
    when 16#0E14# => romdata <= X"FACA455E";
    when 16#0E15# => romdata <= X"6AF96600";
    when 16#0E16# => romdata <= X"AC6FF809";
    when 16#0E17# => romdata <= X"788700DD";
    when 16#0E18# => romdata <= X"2AB93DD2";
    when 16#0E19# => romdata <= X"28483759";
    when 16#0E1A# => romdata <= X"BD903EC0";
    when 16#0E1B# => romdata <= X"02D4C127";
    when 16#0E1C# => romdata <= X"8808B764";
    when 16#0E1D# => romdata <= X"F018E3B7";
    when 16#0E1E# => romdata <= X"40EFD821";
    when 16#0E1F# => romdata <= X"A61F5BEA";
    when 16#0E20# => romdata <= X"2948A653";
    when 16#0E21# => romdata <= X"041FB31F";
    when 16#0E22# => romdata <= X"6D5D0DE0";
    when 16#0E23# => romdata <= X"A045DA36";
    when 16#0E24# => romdata <= X"6E44112C";
    when 16#0E25# => romdata <= X"820FD7FA";
    when 16#0E26# => romdata <= X"966B2CCF";
    when 16#0E27# => romdata <= X"D5A6816A";
    when 16#0E28# => romdata <= X"F84DC0A3";
    when 16#0E29# => romdata <= X"EEB8F9D2";
    when 16#0E2A# => romdata <= X"F0A91258";
    when 16#0E2B# => romdata <= X"6F91D50B";
    when 16#0E2C# => romdata <= X"1AE3D930";
    when 16#0E2D# => romdata <= X"A680A8FB";
    when 16#0E2E# => romdata <= X"7435B687";
    when 16#0E2F# => romdata <= X"5ED2E599";
    when 16#0E30# => romdata <= X"B87598A7";
    when 16#0E31# => romdata <= X"C2024529";
    when 16#0E32# => romdata <= X"6C4965E2";
    when 16#0E33# => romdata <= X"E0CF372B";
    when 16#0E34# => romdata <= X"6ED1219B";
    when 16#0E35# => romdata <= X"A68CB646";
    when 16#0E36# => romdata <= X"D3E73D52";
    when 16#0E37# => romdata <= X"665AAF2E";
    when 16#0E38# => romdata <= X"3D1C4DE8";
    when 16#0E39# => romdata <= X"D2645782";
    when 16#0E3A# => romdata <= X"99B166FA";
    when 16#0E3B# => romdata <= X"0E148281";
    when 16#0E3C# => romdata <= X"C877FA9B";
    when 16#0E3D# => romdata <= X"14818759";
    when 16#0E3E# => romdata <= X"CBF7FF57";
    when 16#0E3F# => romdata <= X"5307E80B";
    when 16#0E40# => romdata <= X"73933599";
    when 16#0E41# => romdata <= X"D94EAD2F";
    when 16#0E42# => romdata <= X"B1C08A30";
    when 16#0E43# => romdata <= X"006330BF";
    when 16#0E44# => romdata <= X"0AC1F1C0";
    when 16#0E45# => romdata <= X"A4EE6B07";
    when 16#0E46# => romdata <= X"F9F3381A";
    when 16#0E47# => romdata <= X"D7E2E469";
    when 16#0E48# => romdata <= X"E8DA9C2D";
    when 16#0E49# => romdata <= X"22CFC0A2";
    when 16#0E4A# => romdata <= X"08B58924";
    when 16#0E4B# => romdata <= X"D2F994AF";
    when 16#0E4C# => romdata <= X"C0268EFE";
    when 16#0E4D# => romdata <= X"206E0A9E";
    when 16#0E4E# => romdata <= X"B79BB51C";
    when 16#0E4F# => romdata <= X"A26FB490";
    when 16#0E50# => romdata <= X"13B9A170";
    when 16#0E51# => romdata <= X"17E0C08F";
    when 16#0E52# => romdata <= X"9FFC6C31";
    when 16#0E53# => romdata <= X"9BB1B5AE";
    when 16#0E54# => romdata <= X"41771443";
    when 16#0E55# => romdata <= X"BC670EEB";
    when 16#0E56# => romdata <= X"91D7769F";
    when 16#0E57# => romdata <= X"9890A9B8";
    when 16#0E58# => romdata <= X"0F52CB01";
    when 16#0E59# => romdata <= X"67EAAF85";
    when 16#0E5A# => romdata <= X"0FAF2A52";
    when 16#0E5B# => romdata <= X"B74ABB17";
    when 16#0E5C# => romdata <= X"92E7CEFF";
    when 16#0E5D# => romdata <= X"68C0D38B";
    when 16#0E5E# => romdata <= X"01F244AC";
    when 16#0E5F# => romdata <= X"0CC0EF07";
    when 16#0E60# => romdata <= X"31E3BDDC";
    when 16#0E61# => romdata <= X"DAB89DF3";
    when 16#0E62# => romdata <= X"76973A7E";
    when 16#0E63# => romdata <= X"D5D4264E";
    when 16#0E64# => romdata <= X"E82C3346";
    when 16#0E65# => romdata <= X"71FCD39E";
    when 16#0E66# => romdata <= X"CD6E2CF8";
    when 16#0E67# => romdata <= X"69493914";
    when 16#0E68# => romdata <= X"F332767B";
    when 16#0E69# => romdata <= X"BE461707";
    when 16#0E6A# => romdata <= X"166A9164";
    when 16#0E6B# => romdata <= X"776D29F5";
    when 16#0E6C# => romdata <= X"EC9291F5";
    when 16#0E6D# => romdata <= X"05AF2912";
    when 16#0E6E# => romdata <= X"54D7319A";
    when 16#0E6F# => romdata <= X"A594B5F3";
    when 16#0E70# => romdata <= X"97D5BDF0";
    when 16#0E71# => romdata <= X"0BB840C4";
    when 16#0E72# => romdata <= X"DDCB425F";
    when 16#0E73# => romdata <= X"4325ED8A";
    when 16#0E74# => romdata <= X"B77E57BE";
    when 16#0E75# => romdata <= X"CA3441B8";
    when 16#0E76# => romdata <= X"94146166";
    when 16#0E77# => romdata <= X"71692EA8";
    when 16#0E78# => romdata <= X"8A89D269";
    when 16#0E79# => romdata <= X"0A4B5FE9";
    when 16#0E7A# => romdata <= X"58F990BD";
    when 16#0E7B# => romdata <= X"84A3884A";
    when 16#0E7C# => romdata <= X"60FADD5D";
    when 16#0E7D# => romdata <= X"A57EDF01";
    when 16#0E7E# => romdata <= X"865F8582";
    when 16#0E7F# => romdata <= X"91954600";
    when 16#0E80# => romdata <= X"B85B6E75";
    when 16#0E81# => romdata <= X"4CC8F680";
    when 16#0E82# => romdata <= X"5A8A19DA";
    when 16#0E83# => romdata <= X"104418D9";
    when 16#0E84# => romdata <= X"C134C8B0";
    when 16#0E85# => romdata <= X"DBCFD5DA";
    when 16#0E86# => romdata <= X"AF5A71BC";
    when 16#0E87# => romdata <= X"047A73BE";
    when 16#0E88# => romdata <= X"DBC192A4";
    when 16#0E89# => romdata <= X"53674BC6";
    when 16#0E8A# => romdata <= X"24959BB7";
    when 16#0E8B# => romdata <= X"6E44C5B3";
    when 16#0E8C# => romdata <= X"4244D473";
    when 16#0E8D# => romdata <= X"6ED3F0F3";
    when 16#0E8E# => romdata <= X"C9658FEC";
    when 16#0E8F# => romdata <= X"0DA5437E";
    when 16#0E90# => romdata <= X"01E12879";
    when 16#0E91# => romdata <= X"5EDD7593";
    when 16#0E92# => romdata <= X"D636CD73";
    when 16#0E93# => romdata <= X"FC1780B3";
    when 16#0E94# => romdata <= X"7A381502";
    when 16#0E95# => romdata <= X"633CCF2E";
    when 16#0E96# => romdata <= X"FDA0BBB4";
    when 16#0E97# => romdata <= X"94C1D0FC";
    when 16#0E98# => romdata <= X"7F602DF8";
    when 16#0E99# => romdata <= X"C282F55E";
    when 16#0E9A# => romdata <= X"3828E81A";
    when 16#0E9B# => romdata <= X"92458EB1";
    when 16#0E9C# => romdata <= X"6B748350";
    when 16#0E9D# => romdata <= X"40D8A9C8";
    when 16#0E9E# => romdata <= X"F2DDF180";
    when 16#0E9F# => romdata <= X"A617B059";
    when 16#0EA0# => romdata <= X"2344B437";
    when 16#0EA1# => romdata <= X"3E1B526C";
    when 16#0EA2# => romdata <= X"9706B843";
    when 16#0EA3# => romdata <= X"B0CED4D2";
    when 16#0EA4# => romdata <= X"5D7324C6";
    when 16#0EA5# => romdata <= X"FDD0F331";
    when 16#0EA6# => romdata <= X"33C00443";
    when 16#0EA7# => romdata <= X"638E6249";
    when 16#0EA8# => romdata <= X"061C56A1";
    when 16#0EA9# => romdata <= X"16CEC782";
    when 16#0EAA# => romdata <= X"2F4512AF";
    when 16#0EAB# => romdata <= X"AEE52CE8";
    when 16#0EAC# => romdata <= X"F94D8547";
    when 16#0EAD# => romdata <= X"F72612EA";
    when 16#0EAE# => romdata <= X"8C7D160C";
    when 16#0EAF# => romdata <= X"65FA3BCC";
    when 16#0EB0# => romdata <= X"92BE0149";
    when 16#0EB1# => romdata <= X"3706EC4E";
    when 16#0EB2# => romdata <= X"5F203F0B";
    when 16#0EB3# => romdata <= X"F85C52F4";
    when 16#0EB4# => romdata <= X"17BAF8AF";
    when 16#0EB5# => romdata <= X"490E5013";
    when 16#0EB6# => romdata <= X"3505685C";
    when 16#0EB7# => romdata <= X"E63AC5B1";
    when 16#0EB8# => romdata <= X"73E07D8D";
    when 16#0EB9# => romdata <= X"ABB2D439";
    when 16#0EBA# => romdata <= X"C6DC18B4";
    when 16#0EBB# => romdata <= X"1B9CF37D";
    when 16#0EBC# => romdata <= X"02C92AB5";
    when 16#0EBD# => romdata <= X"C2F27EC8";
    when 16#0EBE# => romdata <= X"3AB6B2DD";
    when 16#0EBF# => romdata <= X"CB7ABCEA";
    when 16#0EC0# => romdata <= X"30A95BBC";
    when 16#0EC1# => romdata <= X"39E9FD0C";
    when 16#0EC2# => romdata <= X"BB281188";
    when 16#0EC3# => romdata <= X"23F7D034";
    when 16#0EC4# => romdata <= X"2F1EB7B4";
    when 16#0EC5# => romdata <= X"5FA6BB3A";
    when 16#0EC6# => romdata <= X"50223D0D";
    when 16#0EC7# => romdata <= X"7B14E975";
    when 16#0EC8# => romdata <= X"E7658352";
    when 16#0EC9# => romdata <= X"BC9288B4";
    when 16#0ECA# => romdata <= X"8AF13469";
    when 16#0ECB# => romdata <= X"55F4551F";
    when 16#0ECC# => romdata <= X"2ECA47D4";
    when 16#0ECD# => romdata <= X"23EFC63D";
    when 16#0ECE# => romdata <= X"20681057";
    when 16#0ECF# => romdata <= X"E5EF234D";
    when 16#0ED0# => romdata <= X"061A5E6E";
    when 16#0ED1# => romdata <= X"234ED01F";
    when 16#0ED2# => romdata <= X"3DF223A0";
    when 16#0ED3# => romdata <= X"E8B4DEDD";
    when 16#0ED4# => romdata <= X"C552C7DC";
    when 16#0ED5# => romdata <= X"3ECF663D";
    when 16#0ED6# => romdata <= X"5011FC90";
    when 16#0ED7# => romdata <= X"7EB4A7CF";
    when 16#0ED8# => romdata <= X"746AB9E0";
    when 16#0ED9# => romdata <= X"7C2929B7";
    when 16#0EDA# => romdata <= X"427DFE9E";
    when 16#0EDB# => romdata <= X"00B0A130";
    when 16#0EDC# => romdata <= X"88819126";
    when 16#0EDD# => romdata <= X"35A72EA9";
    when 16#0EDE# => romdata <= X"9927F343";
    when 16#0EDF# => romdata <= X"EBAD3243";
    when 16#0EE0# => romdata <= X"6A9B8EB1";
    when 16#0EE1# => romdata <= X"934AC29E";
    when 16#0EE2# => romdata <= X"79BB80AB";
    when 16#0EE3# => romdata <= X"3ED9F5CE";
    when 16#0EE4# => romdata <= X"39D1E43C";
    when 16#0EE5# => romdata <= X"25156465";
    when 16#0EE6# => romdata <= X"4365DA43";
    when 16#0EE7# => romdata <= X"FB8A0FBA";
    when 16#0EE8# => romdata <= X"27F2328D";
    when 16#0EE9# => romdata <= X"82445A1E";
    when 16#0EEA# => romdata <= X"AAED67B9";
    when 16#0EEB# => romdata <= X"2716147E";
    when 16#0EEC# => romdata <= X"859064AC";
    when 16#0EED# => romdata <= X"326A42DC";
    when 16#0EEE# => romdata <= X"7880DE82";
    when 16#0EEF# => romdata <= X"FA782AFF";
    when 16#0EF0# => romdata <= X"F9C59FBD";
    when 16#0EF1# => romdata <= X"CE088746";
    when 16#0EF2# => romdata <= X"F8CEDBA2";
    when 16#0EF3# => romdata <= X"88BC8C2C";
    when 16#0EF4# => romdata <= X"4B458782";
    when 16#0EF5# => romdata <= X"CC9BE63A";
    when 16#0EF6# => romdata <= X"86168B67";
    when 16#0EF7# => romdata <= X"1BE99A09";
    when 16#0EF8# => romdata <= X"F2217B7B";
    when 16#0EF9# => romdata <= X"B2A7BC88";
    when 16#0EFA# => romdata <= X"651C1BCE";
    when 16#0EFB# => romdata <= X"8A0B8931";
    when 16#0EFC# => romdata <= X"6ABFE72B";
    when 16#0EFD# => romdata <= X"22722273";
    when 16#0EFE# => romdata <= X"AF570974";
    when 16#0EFF# => romdata <= X"D8EDEE40";
    when 16#0F00# => romdata <= X"DD40DD43";
    when 16#0F01# => romdata <= X"8251E401";
    when 16#0F02# => romdata <= X"FC926CC6";
    when 16#0F03# => romdata <= X"96839341";
    when 16#0F04# => romdata <= X"5D52D521";
    when 16#0F05# => romdata <= X"A5BB34D4";
    when 16#0F06# => romdata <= X"272D6BC7";
    when 16#0F07# => romdata <= X"B5431062";
    when 16#0F08# => romdata <= X"B35112CA";
    when 16#0F09# => romdata <= X"709C0680";
    when 16#0F0A# => romdata <= X"CBB18EEE";
    when 16#0F0B# => romdata <= X"053AAD62";
    when 16#0F0C# => romdata <= X"B2391C9E";
    when 16#0F0D# => romdata <= X"9D580562";
    when 16#0F0E# => romdata <= X"541A453E";
    when 16#0F0F# => romdata <= X"D936CE8E";
    when 16#0F10# => romdata <= X"88DFA61A";
    when 16#0F11# => romdata <= X"88CA3BEE";
    when 16#0F12# => romdata <= X"66CFFF80";
    when 16#0F13# => romdata <= X"1785CCE8";
    when 16#0F14# => romdata <= X"63ED9C36";
    when 16#0F15# => romdata <= X"A04D2DC8";
    when 16#0F16# => romdata <= X"742A81CA";
    when 16#0F17# => romdata <= X"55127B44";
    when 16#0F18# => romdata <= X"314AB4E6";
    when 16#0F19# => romdata <= X"87ED921B";
    when 16#0F1A# => romdata <= X"4881CB36";
    when 16#0F1B# => romdata <= X"3AFB3CCE";
    when 16#0F1C# => romdata <= X"7EB774E3";
    when 16#0F1D# => romdata <= X"205D4591";
    when 16#0F1E# => romdata <= X"939ED7D3";
    when 16#0F1F# => romdata <= X"C0C508A3";
    when 16#0F20# => romdata <= X"1786421F";
    when 16#0F21# => romdata <= X"49669E12";
    when 16#0F22# => romdata <= X"0F01D35D";
    when 16#0F23# => romdata <= X"467B40F8";
    when 16#0F24# => romdata <= X"5F2454F1";
    when 16#0F25# => romdata <= X"3F591F3B";
    when 16#0F26# => romdata <= X"83093742";
    when 16#0F27# => romdata <= X"1B5C8A6C";
    when 16#0F28# => romdata <= X"20EA8789";
    when 16#0F29# => romdata <= X"71AEC941";
    when 16#0F2A# => romdata <= X"FD99CEA9";
    when 16#0F2B# => romdata <= X"2FEE00E5";
    when 16#0F2C# => romdata <= X"DC226498";
    when 16#0F2D# => romdata <= X"7DBC549E";
    when 16#0F2E# => romdata <= X"FF3E4A26";
    when 16#0F2F# => romdata <= X"AF0CAD74";
    when 16#0F30# => romdata <= X"21C4256D";
    when 16#0F31# => romdata <= X"107A3E89";
    when 16#0F32# => romdata <= X"08F67450";
    when 16#0F33# => romdata <= X"960E4E41";
    when 16#0F34# => romdata <= X"FD7E2E84";
    when 16#0F35# => romdata <= X"F754BAC8";
    when 16#0F36# => romdata <= X"1C8F5F1D";
    when 16#0F37# => romdata <= X"6F650DEB";
    when 16#0F38# => romdata <= X"3E6EFF60";
    when 16#0F39# => romdata <= X"59836643";
    when 16#0F3A# => romdata <= X"209E3880";
    when 16#0F3B# => romdata <= X"D7BDA701";
    when 16#0F3C# => romdata <= X"869208D8";
    when 16#0F3D# => romdata <= X"E4BC8D06";
    when 16#0F3E# => romdata <= X"14066414";
    when 16#0F3F# => romdata <= X"DB3F93D6";
    when 16#0F40# => romdata <= X"EA187950";
    when 16#0F41# => romdata <= X"285F55BB";
    when 16#0F42# => romdata <= X"7A1B026E";
    when 16#0F43# => romdata <= X"A4BFCAB4";
    when 16#0F44# => romdata <= X"671B0770";
    when 16#0F45# => romdata <= X"4828D5CB";
    when 16#0F46# => romdata <= X"F9730EFC";
    when 16#0F47# => romdata <= X"99E68E91";
    when 16#0F48# => romdata <= X"F1FE9664";
    when 16#0F49# => romdata <= X"DFA73297";
    when 16#0F4A# => romdata <= X"F2D6BD94";
    when 16#0F4B# => romdata <= X"97DE0498";
    when 16#0F4C# => romdata <= X"2C9FF373";
    when 16#0F4D# => romdata <= X"0BB6FC3E";
    when 16#0F4E# => romdata <= X"A2053B3F";
    when 16#0F4F# => romdata <= X"45DC7FB5";
    when 16#0F50# => romdata <= X"87BA19B3";
    when 16#0F51# => romdata <= X"C6B7E780";
    when 16#0F52# => romdata <= X"EA5F25B4";
    when 16#0F53# => romdata <= X"5BB72717";
    when 16#0F54# => romdata <= X"4D4CD3B4";
    when 16#0F55# => romdata <= X"01FE1906";
    when 16#0F56# => romdata <= X"360BF0B1";
    when 16#0F57# => romdata <= X"5DB13B62";
    when 16#0F58# => romdata <= X"752F82EC";
    when 16#0F59# => romdata <= X"62226AAB";
    when 16#0F5A# => romdata <= X"C83C1C26";
    when 16#0F5B# => romdata <= X"376F8366";
    when 16#0F5C# => romdata <= X"BB849DDB";
    when 16#0F5D# => romdata <= X"65958AD9";
    when 16#0F5E# => romdata <= X"69B25654";
    when 16#0F5F# => romdata <= X"DEF18415";
    when 16#0F60# => romdata <= X"18993033";
    when 16#0F61# => romdata <= X"AF47EABE";
    when 16#0F62# => romdata <= X"E3CAAA93";
    when 16#0F63# => romdata <= X"6F19E28A";
    when 16#0F64# => romdata <= X"205F3CDD";
    when 16#0F65# => romdata <= X"B5CAC649";
    when 16#0F66# => romdata <= X"DB6A9048";
    when 16#0F67# => romdata <= X"3ACB63A2";
    when 16#0F68# => romdata <= X"4EA46D39";
    when 16#0F69# => romdata <= X"7508EEB5";
    when 16#0F6A# => romdata <= X"DA94E9C8";
    when 16#0F6B# => romdata <= X"83EB0451";
    when 16#0F6C# => romdata <= X"D036E28C";
    when 16#0F6D# => romdata <= X"C303D52B";
    when 16#0F6E# => romdata <= X"1BB31FFF";
    when 16#0F6F# => romdata <= X"582605F3";
    when 16#0F70# => romdata <= X"40D44950";
    when 16#0F71# => romdata <= X"8959ED1F";
    when 16#0F72# => romdata <= X"E2FF0BD2";
    when 16#0F73# => romdata <= X"2FDF77F9";
    when 16#0F74# => romdata <= X"680D6B56";
    when 16#0F75# => romdata <= X"47D59E7E";
    when 16#0F76# => romdata <= X"6A003AF0";
    when 16#0F77# => romdata <= X"C6A95092";
    when 16#0F78# => romdata <= X"F0DE43D1";
    when 16#0F79# => romdata <= X"252EA6DE";
    when 16#0F7A# => romdata <= X"00F288BC";
    when 16#0F7B# => romdata <= X"CE3ED9CE";
    when 16#0F7C# => romdata <= X"273DCB4F";
    when 16#0F7D# => romdata <= X"3BA7E8D1";
    when 16#0F7E# => romdata <= X"7353B8EC";
    when 16#0F7F# => romdata <= X"A24F03A0";
    when 16#0F80# => romdata <= X"FE38B1AC";
    when 16#0F81# => romdata <= X"A366B4C1";
    when 16#0F82# => romdata <= X"5F3FDD4D";
    when 16#0F83# => romdata <= X"F0E0274F";
    when 16#0F84# => romdata <= X"BEFDA004";
    when 16#0F85# => romdata <= X"2BB203A4";
    when 16#0F86# => romdata <= X"F6627ED9";
    when 16#0F87# => romdata <= X"E29F4053";
    when 16#0F88# => romdata <= X"79B2F2DD";
    when 16#0F89# => romdata <= X"C0F3B02A";
    when 16#0F8A# => romdata <= X"0CA70A94";
    when 16#0F8B# => romdata <= X"99F3CE82";
    when 16#0F8C# => romdata <= X"B87603FA";
    when 16#0F8D# => romdata <= X"A347B705";
    when 16#0F8E# => romdata <= X"2CB5D13D";
    when 16#0F8F# => romdata <= X"9DE84C11";
    when 16#0F90# => romdata <= X"4EF3B8F6";
    when 16#0F91# => romdata <= X"2418FB1F";
    when 16#0F92# => romdata <= X"3E374B99";
    when 16#0F93# => romdata <= X"7127667F";
    when 16#0F94# => romdata <= X"D6BCA2E2";
    when 16#0F95# => romdata <= X"F9DBC04E";
    when 16#0F96# => romdata <= X"CA9D908C";
    when 16#0F97# => romdata <= X"D37C62F0";
    when 16#0F98# => romdata <= X"8EEA6F44";
    when 16#0F99# => romdata <= X"B3FDC149";
    when 16#0F9A# => romdata <= X"465AA803";
    when 16#0F9B# => romdata <= X"7D65A6C8";
    when 16#0F9C# => romdata <= X"B9B8B3D5";
    when 16#0F9D# => romdata <= X"E9A40578";
    when 16#0F9E# => romdata <= X"E5EA3AE1";
    when 16#0F9F# => romdata <= X"209BA49E";
    when 16#0FA0# => romdata <= X"5E2AC615";
    when 16#0FA1# => romdata <= X"C59A2D71";
    when 16#0FA2# => romdata <= X"AC1605B9";
    when 16#0FA3# => romdata <= X"8E39A5E6";
    when 16#0FA4# => romdata <= X"6A890754";
    when 16#0FA5# => romdata <= X"C7D1C07E";
    when 16#0FA6# => romdata <= X"06DE7863";
    when 16#0FA7# => romdata <= X"2587BADA";
    when 16#0FA8# => romdata <= X"F7FAAB0A";
    when 16#0FA9# => romdata <= X"529AB791";
    when 16#0FAA# => romdata <= X"095DB0A7";
    when 16#0FAB# => romdata <= X"08B691E9";
    when 16#0FAC# => romdata <= X"D81F2CEA";
    when 16#0FAD# => romdata <= X"8F07B054";
    when 16#0FAE# => romdata <= X"95528B9F";
    when 16#0FAF# => romdata <= X"D56F77A4";
    when 16#0FB0# => romdata <= X"C8209DB9";
    when 16#0FB1# => romdata <= X"72FAADD9";
    when 16#0FB2# => romdata <= X"791BA59F";
    when 16#0FB3# => romdata <= X"47C06F24";
    when 16#0FB4# => romdata <= X"1F50C061";
    when 16#0FB5# => romdata <= X"9FC04F84";
    when 16#0FB6# => romdata <= X"56339E0A";
    when 16#0FB7# => romdata <= X"F331310F";
    when 16#0FB8# => romdata <= X"A4DCCBEA";
    when 16#0FB9# => romdata <= X"0E5DC279";
    when 16#0FBA# => romdata <= X"5CA6B3AD";
    when 16#0FBB# => romdata <= X"D0174AE4";
    when 16#0FBC# => romdata <= X"B30AC042";
    when 16#0FBD# => romdata <= X"8320ACEA";
    when 16#0FBE# => romdata <= X"FF68F73E";
    when 16#0FBF# => romdata <= X"D11DC1BC";
    when 16#0FC0# => romdata <= X"9F0237BD";
    when 16#0FC1# => romdata <= X"C75F7F48";
    when 16#0FC2# => romdata <= X"BE518EB3";
    when 16#0FC3# => romdata <= X"305CF2BB";
    when 16#0FC4# => romdata <= X"898B3297";
    when 16#0FC5# => romdata <= X"16FC9ECF";
    when 16#0FC6# => romdata <= X"7E99B510";
    when 16#0FC7# => romdata <= X"B3309808";
    when 16#0FC8# => romdata <= X"735FD0A7";
    when 16#0FC9# => romdata <= X"7B15731C";
    when 16#0FCA# => romdata <= X"233998F9";
    when 16#0FCB# => romdata <= X"ECEF46E2";
    when 16#0FCC# => romdata <= X"CAA6E6ED";
    when 16#0FCD# => romdata <= X"C8D05B94";
    when 16#0FCE# => romdata <= X"3ABD1702";
    when 16#0FCF# => romdata <= X"7A80D636";
    when 16#0FD0# => romdata <= X"E535038F";
    when 16#0FD1# => romdata <= X"AE44D60A";
    when 16#0FD2# => romdata <= X"AEC5406A";
    when 16#0FD3# => romdata <= X"372D6247";
    when 16#0FD4# => romdata <= X"9192FA84";
    when 16#0FD5# => romdata <= X"D844520C";
    when 16#0FD6# => romdata <= X"6774CC58";
    when 16#0FD7# => romdata <= X"9FEE16A3";
    when 16#0FD8# => romdata <= X"A5549495";
    when 16#0FD9# => romdata <= X"D968AABA";
    when 16#0FDA# => romdata <= X"ABFE4DB9";
    when 16#0FDB# => romdata <= X"4F5AE0C5";
    when 16#0FDC# => romdata <= X"4E603D6D";
    when 16#0FDD# => romdata <= X"A5C30567";
    when 16#0FDE# => romdata <= X"69A06489";
    when 16#0FDF# => romdata <= X"0533EA8E";
    when 16#0FE0# => romdata <= X"A1E5D1CD";
    when 16#0FE1# => romdata <= X"410CC8DD";
    when 16#0FE2# => romdata <= X"4B1D7E0F";
    when 16#0FE3# => romdata <= X"5F787232";
    when 16#0FE4# => romdata <= X"439AA4B3";
    when 16#0FE5# => romdata <= X"911C5DC7";
    when 16#0FE6# => romdata <= X"92ECB873";
    when 16#0FE7# => romdata <= X"E8105A1A";
    when 16#0FE8# => romdata <= X"A61C627B";
    when 16#0FE9# => romdata <= X"E57E809C";
    when 16#0FEA# => romdata <= X"6863073E";
    when 16#0FEB# => romdata <= X"1E19AD8B";
    when 16#0FEC# => romdata <= X"987DE97D";
    when 16#0FED# => romdata <= X"88A817FB";
    when 16#0FEE# => romdata <= X"43ADBB77";
    when 16#0FEF# => romdata <= X"51E36D1F";
    when 16#0FF0# => romdata <= X"0E7B70B3";
    when 16#0FF1# => romdata <= X"759D6EA8";
    when 16#0FF2# => romdata <= X"F2350D10";
    when 16#0FF3# => romdata <= X"AF38C331";
    when 16#0FF4# => romdata <= X"E22703B2";
    when 16#0FF5# => romdata <= X"B5103C90";
    when 16#0FF6# => romdata <= X"8E1D35A8";
    when 16#0FF7# => romdata <= X"E814E45B";
    when 16#0FF8# => romdata <= X"AE81DCA0";
    when 16#0FF9# => romdata <= X"530FC352";
    when 16#0FFA# => romdata <= X"5CD64054";
    when 16#0FFB# => romdata <= X"8245C259";
    when 16#0FFC# => romdata <= X"738E749E";
    when 16#0FFD# => romdata <= X"195B0060";
    when 16#0FFE# => romdata <= X"81A18C45";
    when 16#0FFF# => romdata <= X"475F9060";
    when 16#1000# => romdata <= X"B39340CA";
    when 16#1001# => romdata <= X"1C817D81";
    when 16#1002# => romdata <= X"EF4FAE4E";
    when 16#1003# => romdata <= X"95BF3504";
    when 16#1004# => romdata <= X"A7709089";
    when 16#1005# => romdata <= X"FB48560E";
    when 16#1006# => romdata <= X"9E3EF802";
    when 16#1007# => romdata <= X"180E85EB";
    when 16#1008# => romdata <= X"2194E059";
    when 16#1009# => romdata <= X"02C6C4C5";
    when 16#100A# => romdata <= X"2021FEB7";
    when 16#100B# => romdata <= X"EC64FD41";
    when 16#100C# => romdata <= X"6BCEBC8E";
    when 16#100D# => romdata <= X"39D64A4B";
    when 16#100E# => romdata <= X"5EE34529";
    when 16#100F# => romdata <= X"1911AB82";
    when 16#1010# => romdata <= X"04A888C2";
    when 16#1011# => romdata <= X"5B1CD3D9";
    when 16#1012# => romdata <= X"342A56C5";
    when 16#1013# => romdata <= X"38636D3E";
    when 16#1014# => romdata <= X"AB957037";
    when 16#1015# => romdata <= X"D09E879A";
    when 16#1016# => romdata <= X"E5F3A398";
    when 16#1017# => romdata <= X"34FBB84A";
    when 16#1018# => romdata <= X"3D8D5090";
    when 16#1019# => romdata <= X"D7814246";
    when 16#101A# => romdata <= X"B62E9CA6";
    when 16#101B# => romdata <= X"8533D2EC";
    when 16#101C# => romdata <= X"403B4FB9";
    when 16#101D# => romdata <= X"488467FF";
    when 16#101E# => romdata <= X"9758B0D1";
    when 16#101F# => romdata <= X"5A8CEF89";
    when 16#1020# => romdata <= X"187A1D58";
    when 16#1021# => romdata <= X"97880040";
    when 16#1022# => romdata <= X"B6C3C524";
    when 16#1023# => romdata <= X"4E85A2AD";
    when 16#1024# => romdata <= X"14BCF2F5";
    when 16#1025# => romdata <= X"ABC44A7B";
    when 16#1026# => romdata <= X"1D4A87E8";
    when 16#1027# => romdata <= X"BDA05766";
    when 16#1028# => romdata <= X"218773ED";
    when 16#1029# => romdata <= X"4F70F8D1";
    when 16#102A# => romdata <= X"D07CBB1E";
    when 16#102B# => romdata <= X"8CA6298E";
    when 16#102C# => romdata <= X"64EE6DC5";
    when 16#102D# => romdata <= X"886D3749";
    when 16#102E# => romdata <= X"5BA2EDB3";
    when 16#102F# => romdata <= X"E0B0B68A";
    when 16#1030# => romdata <= X"D9F30031";
    when 16#1031# => romdata <= X"0B88898D";
    when 16#1032# => romdata <= X"DEEFD484";
    when 16#1033# => romdata <= X"538C31A9";
    when 16#1034# => romdata <= X"BCAA76EC";
    when 16#1035# => romdata <= X"AD0C1660";
    when 16#1036# => romdata <= X"7D321890";
    when 16#1037# => romdata <= X"58B0862E";
    when 16#1038# => romdata <= X"E9D70CEA";
    when 16#1039# => romdata <= X"9D304755";
    when 16#103A# => romdata <= X"CE8037BA";
    when 16#103B# => romdata <= X"4C46C257";
    when 16#103C# => romdata <= X"3181748A";
    when 16#103D# => romdata <= X"212E4B2B";
    when 16#103E# => romdata <= X"DD04F9BC";
    when 16#103F# => romdata <= X"24051827";
    when 16#1040# => romdata <= X"3DC17CBA";
    when 16#1041# => romdata <= X"FF21A03E";
    when 16#1042# => romdata <= X"9120FA7D";
    when 16#1043# => romdata <= X"CA18D56D";
    when 16#1044# => romdata <= X"D1D9A7E5";
    when 16#1045# => romdata <= X"10C90CF2";
    when 16#1046# => romdata <= X"19104385";
    when 16#1047# => romdata <= X"F531F2EF";
    when 16#1048# => romdata <= X"AFD185EC";
    when 16#1049# => romdata <= X"B6B911F9";
    when 16#104A# => romdata <= X"B7809D98";
    when 16#104B# => romdata <= X"D86F1551";
    when 16#104C# => romdata <= X"6FFDDBE9";
    when 16#104D# => romdata <= X"BD1CF866";
    when 16#104E# => romdata <= X"2EB777C3";
    when 16#104F# => romdata <= X"F94EA3F9";
    when 16#1050# => romdata <= X"62D7B794";
    when 16#1051# => romdata <= X"49FAAD39";
    when 16#1052# => romdata <= X"935429E9";
    when 16#1053# => romdata <= X"2CAE5637";
    when 16#1054# => romdata <= X"E9BCF4E9";
    when 16#1055# => romdata <= X"4D413D27";
    when 16#1056# => romdata <= X"93495240";
    when 16#1057# => romdata <= X"9AB536BE";
    when 16#1058# => romdata <= X"4055AFBC";
    when 16#1059# => romdata <= X"4330CD1E";
    when 16#105A# => romdata <= X"4B5509EF";
    when 16#105B# => romdata <= X"E5F8EFC9";
    when 16#105C# => romdata <= X"ECBE9EF3";
    when 16#105D# => romdata <= X"77DE7E37";
    when 16#105E# => romdata <= X"C479BB9D";
    when 16#105F# => romdata <= X"3EE7745E";
    when 16#1060# => romdata <= X"4609B0A6";
    when 16#1061# => romdata <= X"D2C5D92E";
    when 16#1062# => romdata <= X"B3C9E227";
    when 16#1063# => romdata <= X"8C1F2221";
    when 16#1064# => romdata <= X"FF907596";
    when 16#1065# => romdata <= X"AA5E096A";
    when 16#1066# => romdata <= X"CF8990EB";
    when 16#1067# => romdata <= X"A907E43A";
    when 16#1068# => romdata <= X"D320F801";
    when 16#1069# => romdata <= X"9CB6355A";
    when 16#106A# => romdata <= X"2BA8670E";
    when 16#106B# => romdata <= X"E5A4F463";
    when 16#106C# => romdata <= X"E8E56F8F";
    when 16#106D# => romdata <= X"1D3E7F49";
    when 16#106E# => romdata <= X"22510FB6";
    when 16#106F# => romdata <= X"68E32C4C";
    when 16#1070# => romdata <= X"F23AD849";
    when 16#1071# => romdata <= X"6399638B";
    when 16#1072# => romdata <= X"095B4783";
    when 16#1073# => romdata <= X"3E0CBB34";
    when 16#1074# => romdata <= X"977EB3E4";
    when 16#1075# => romdata <= X"242EAF87";
    when 16#1076# => romdata <= X"0D86660D";
    when 16#1077# => romdata <= X"6A73F83E";
    when 16#1078# => romdata <= X"45D6E8A4";
    when 16#1079# => romdata <= X"1EDCA381";
    when 16#107A# => romdata <= X"50796495";
    when 16#107B# => romdata <= X"44597C5C";
    when 16#107C# => romdata <= X"43B6C93F";
    when 16#107D# => romdata <= X"EBAD5700";
    when 16#107E# => romdata <= X"D22EDAF4";
    when 16#107F# => romdata <= X"31FD3400";
    when 16#1080# => romdata <= X"A64F94BB";
    when 16#1081# => romdata <= X"47BD4033";
    when 16#1082# => romdata <= X"C76D4924";
    when 16#1083# => romdata <= X"305907EC";
    when 16#1084# => romdata <= X"1F618B43";
    when 16#1085# => romdata <= X"C7535F3C";
    when 16#1086# => romdata <= X"FC093E5A";
    when 16#1087# => romdata <= X"F5DDD5C4";
    when 16#1088# => romdata <= X"339F3BB6";
    when 16#1089# => romdata <= X"D835B5C2";
    when 16#108A# => romdata <= X"C2053CD3";
    when 16#108B# => romdata <= X"D5693368";
    when 16#108C# => romdata <= X"D4E1A7CA";
    when 16#108D# => romdata <= X"C59425D1";
    when 16#108E# => romdata <= X"FD96809C";
    when 16#108F# => romdata <= X"67285CFD";
    when 16#1090# => romdata <= X"3FC05B01";
    when 16#1091# => romdata <= X"053CB077";
    when 16#1092# => romdata <= X"3221D720";
    when 16#1093# => romdata <= X"5778022F";
    when 16#1094# => romdata <= X"487BF99D";
    when 16#1095# => romdata <= X"1650566B";
    when 16#1096# => romdata <= X"E287FD7A";
    when 16#1097# => romdata <= X"E882AA8E";
    when 16#1098# => romdata <= X"8F52E5D4";
    when 16#1099# => romdata <= X"E3C0C2F9";
    when 16#109A# => romdata <= X"71C9FF70";
    when 16#109B# => romdata <= X"AA378691";
    when 16#109C# => romdata <= X"EBD8ADE4";
    when 16#109D# => romdata <= X"5CF21382";
    when 16#109E# => romdata <= X"2D09FD05";
    when 16#109F# => romdata <= X"243F9726";
    when 16#10A0# => romdata <= X"F6C69893";
    when 16#10A1# => romdata <= X"845E57C3";
    when 16#10A2# => romdata <= X"7A7643E1";
    when 16#10A3# => romdata <= X"6B770E26";
    when 16#10A4# => romdata <= X"F431FF69";
    when 16#10A5# => romdata <= X"D4372719";
    when 16#10A6# => romdata <= X"05D270EB";
    when 16#10A7# => romdata <= X"85D8D229";
    when 16#10A8# => romdata <= X"D7D87662";
    when 16#10A9# => romdata <= X"121F0BEE";
    when 16#10AA# => romdata <= X"B1E895ED";
    when 16#10AB# => romdata <= X"9589A9CF";
    when 16#10AC# => romdata <= X"5833408A";
    when 16#10AD# => romdata <= X"04197AC9";
    when 16#10AE# => romdata <= X"025D8570";
    when 16#10AF# => romdata <= X"AD9B75DB";
    when 16#10B0# => romdata <= X"7E192EA0";
    when 16#10B1# => romdata <= X"A0895049";
    when 16#10B2# => romdata <= X"96E9DC65";
    when 16#10B3# => romdata <= X"2975D836";
    when 16#10B4# => romdata <= X"33619CFF";
    when 16#10B5# => romdata <= X"80667D8B";
    when 16#10B6# => romdata <= X"519536B3";
    when 16#10B7# => romdata <= X"475248BA";
    when 16#10B8# => romdata <= X"8213C8A4";
    when 16#10B9# => romdata <= X"C66DE69B";
    when 16#10BA# => romdata <= X"4B3774BF";
    when 16#10BB# => romdata <= X"9142425C";
    when 16#10BC# => romdata <= X"57F34A27";
    when 16#10BD# => romdata <= X"B1E28811";
    when 16#10BE# => romdata <= X"9E3FFCC6";
    when 16#10BF# => romdata <= X"AF6A2108";
    when 16#10C0# => romdata <= X"7F9394F0";
    when 16#10C1# => romdata <= X"9DDFBD42";
    when 16#10C2# => romdata <= X"F32D059B";
    when 16#10C3# => romdata <= X"8CD4104A";
    when 16#10C4# => romdata <= X"519BA640";
    when 16#10C5# => romdata <= X"765D5CDE";
    when 16#10C6# => romdata <= X"490E62F1";
    when 16#10C7# => romdata <= X"0E695FBF";
    when 16#10C8# => romdata <= X"D33CBC9D";
    when 16#10C9# => romdata <= X"2208A532";
    when 16#10CA# => romdata <= X"C8EC25DA";
    when 16#10CB# => romdata <= X"28B8CC1B";
    when 16#10CC# => romdata <= X"6850AB43";
    when 16#10CD# => romdata <= X"D9B5C00B";
    when 16#10CE# => romdata <= X"6E74B7A1";
    when 16#10CF# => romdata <= X"48791AB0";
    when 16#10D0# => romdata <= X"7B328D34";
    when 16#10D1# => romdata <= X"7058C7E6";
    when 16#10D2# => romdata <= X"233E18C5";
    when 16#10D3# => romdata <= X"ED172C9F";
    when 16#10D4# => romdata <= X"9E9ACF29";
    when 16#10D5# => romdata <= X"D913E2A1";
    when 16#10D6# => romdata <= X"614BFC08";
    when 16#10D7# => romdata <= X"93D4967E";
    when 16#10D8# => romdata <= X"D033B2B9";
    when 16#10D9# => romdata <= X"AE6B51F9";
    when 16#10DA# => romdata <= X"08F1CED5";
    when 16#10DB# => romdata <= X"7C14FEEA";
    when 16#10DC# => romdata <= X"85CD4D97";
    when 16#10DD# => romdata <= X"11216BE7";
    when 16#10DE# => romdata <= X"F79FA672";
    when 16#10DF# => romdata <= X"1B7DCCA0";
    when 16#10E0# => romdata <= X"33C80127";
    when 16#10E1# => romdata <= X"AC6E5FCF";
    when 16#10E2# => romdata <= X"58EB4005";
    when 16#10E3# => romdata <= X"EC24CB48";
    when 16#10E4# => romdata <= X"86D78735";
    when 16#10E5# => romdata <= X"5362D5E7";
    when 16#10E6# => romdata <= X"031B9B2A";
    when 16#10E7# => romdata <= X"C2A86D73";
    when 16#10E8# => romdata <= X"0AD73418";
    when 16#10E9# => romdata <= X"1E723A81";
    when 16#10EA# => romdata <= X"1FF510A4";
    when 16#10EB# => romdata <= X"DF868001";
    when 16#10EC# => romdata <= X"973FE832";
    when 16#10ED# => romdata <= X"88D78E6F";
    when 16#10EE# => romdata <= X"9B9441DA";
    when 16#10EF# => romdata <= X"F5BE2974";
    when 16#10F0# => romdata <= X"A2848FD9";
    when 16#10F1# => romdata <= X"17C3BCD3";
    when 16#10F2# => romdata <= X"46A43192";
    when 16#10F3# => romdata <= X"2246EC85";
    when 16#10F4# => romdata <= X"2E4AAD46";
    when 16#10F5# => romdata <= X"7E60C15D";
    when 16#10F6# => romdata <= X"61DD3BF4";
    when 16#10F7# => romdata <= X"A207BB57";
    when 16#10F8# => romdata <= X"DB45DCAD";
    when 16#10F9# => romdata <= X"EFE3210B";
    when 16#10FA# => romdata <= X"E74B9DAC";
    when 16#10FB# => romdata <= X"C918A394";
    when 16#10FC# => romdata <= X"469F2E2C";
    when 16#10FD# => romdata <= X"95AD1E21";
    when 16#10FE# => romdata <= X"1947948F";
    when 16#10FF# => romdata <= X"E24F5E40";
    when 16#1100# => romdata <= X"FD1F6976";
    when 16#1101# => romdata <= X"002C39C8";
    when 16#1102# => romdata <= X"7187C44E";
    when 16#1103# => romdata <= X"3D224ED4";
    when 16#1104# => romdata <= X"DF0B6775";
    when 16#1105# => romdata <= X"0105944C";
    when 16#1106# => romdata <= X"651A5E57";
    when 16#1107# => romdata <= X"798F168A";
    when 16#1108# => romdata <= X"136AC0FB";
    when 16#1109# => romdata <= X"5979C4E8";
    when 16#110A# => romdata <= X"47A82B20";
    when 16#110B# => romdata <= X"A2E6C45D";
    when 16#110C# => romdata <= X"B42EF2B9";
    when 16#110D# => romdata <= X"30A80D32";
    when 16#110E# => romdata <= X"57BCCC53";
    when 16#110F# => romdata <= X"EDA966F5";
    when 16#1110# => romdata <= X"DCD9AD47";
    when 16#1111# => romdata <= X"CFB226EE";
    when 16#1112# => romdata <= X"D9B62A87";
    when 16#1113# => romdata <= X"4E9F6404";
    when 16#1114# => romdata <= X"D4087798";
    when 16#1115# => romdata <= X"A1005F41";
    when 16#1116# => romdata <= X"31171D3A";
    when 16#1117# => romdata <= X"47907A3C";
    when 16#1118# => romdata <= X"D602B83D";
    when 16#1119# => romdata <= X"ABE094D2";
    when 16#111A# => romdata <= X"CB031867";
    when 16#111B# => romdata <= X"DF4595F3";
    when 16#111C# => romdata <= X"ED59FD8C";
    when 16#111D# => romdata <= X"4D76EDEE";
    when 16#111E# => romdata <= X"E59E422C";
    when 16#111F# => romdata <= X"E5C7D0A5";
    when 16#1120# => romdata <= X"F720BE94";
    when 16#1121# => romdata <= X"FA24DF05";
    when 16#1122# => romdata <= X"F758348E";
    when 16#1123# => romdata <= X"ADD5EFE9";
    when 16#1124# => romdata <= X"197C6BB2";
    when 16#1125# => romdata <= X"292E2B14";
    when 16#1126# => romdata <= X"DB8C6DB2";
    when 16#1127# => romdata <= X"4AA94C5F";
    when 16#1128# => romdata <= X"F0F5106D";
    when 16#1129# => romdata <= X"2B566058";
    when 16#112A# => romdata <= X"D32C58B6";
    when 16#112B# => romdata <= X"3A150784";
    when 16#112C# => romdata <= X"F7B02478";
    when 16#112D# => romdata <= X"D9973DD4";
    when 16#112E# => romdata <= X"CFD2E840";
    when 16#112F# => romdata <= X"59AE0F4F";
    when 16#1130# => romdata <= X"1320754B";
    when 16#1131# => romdata <= X"7EE83F04";
    when 16#1132# => romdata <= X"A51C67EF";
    when 16#1133# => romdata <= X"FC2EB1C3";
    when 16#1134# => romdata <= X"01C0C58D";
    when 16#1135# => romdata <= X"BAEBE954";
    when 16#1136# => romdata <= X"74E3484A";
    when 16#1137# => romdata <= X"76500103";
    when 16#1138# => romdata <= X"C14C40BB";
    when 16#1139# => romdata <= X"0B7D3A04";
    when 16#113A# => romdata <= X"D8BDABB6";
    when 16#113B# => romdata <= X"05C1EF9F";
    when 16#113C# => romdata <= X"D4A65649";
    when 16#113D# => romdata <= X"34DEC50B";
    when 16#113E# => romdata <= X"D5878243";
    when 16#113F# => romdata <= X"AEE80F97";
    when 16#1140# => romdata <= X"96EED70C";
    when 16#1141# => romdata <= X"E1B1E8B5";
    when 16#1142# => romdata <= X"5725DF76";
    when 16#1143# => romdata <= X"472D12D4";
    when 16#1144# => romdata <= X"A7A48798";
    when 16#1145# => romdata <= X"9F42E670";
    when 16#1146# => romdata <= X"5818B1F7";
    when 16#1147# => romdata <= X"E149E971";
    when 16#1148# => romdata <= X"53A7B05A";
    when 16#1149# => romdata <= X"82FA3FBE";
    when 16#114A# => romdata <= X"51763E61";
    when 16#114B# => romdata <= X"171A4E12";
    when 16#114C# => romdata <= X"931472E9";
    when 16#114D# => romdata <= X"4CCBA74C";
    when 16#114E# => romdata <= X"C09483DF";
    when 16#114F# => romdata <= X"93623FC6";
    when 16#1150# => romdata <= X"0945070F";
    when 16#1151# => romdata <= X"DDF3A00B";
    when 16#1152# => romdata <= X"56165042";
    when 16#1153# => romdata <= X"7E4BD64D";
    when 16#1154# => romdata <= X"675B1EB3";
    when 16#1155# => romdata <= X"98B35EF0";
    when 16#1156# => romdata <= X"57A66FD0";
    when 16#1157# => romdata <= X"B48EDBAB";
    when 16#1158# => romdata <= X"BDCD57C3";
    when 16#1159# => romdata <= X"2ABAE46F";
    when 16#115A# => romdata <= X"5CDD0CB1";
    when 16#115B# => romdata <= X"FCF17765";
    when 16#115C# => romdata <= X"258236F3";
    when 16#115D# => romdata <= X"DE40BD5D";
    when 16#115E# => romdata <= X"0A3C5C97";
    when 16#115F# => romdata <= X"8D81DEB0";
    when 16#1160# => romdata <= X"7367AB20";
    when 16#1161# => romdata <= X"B2CAA983";
    when 16#1162# => romdata <= X"4B957616";
    when 16#1163# => romdata <= X"1C4F20FB";
    when 16#1164# => romdata <= X"9C184A01";
    when 16#1165# => romdata <= X"DC9021A4";
    when 16#1166# => romdata <= X"E92B7133";
    when 16#1167# => romdata <= X"3354E05B";
    when 16#1168# => romdata <= X"BEA9015E";
    when 16#1169# => romdata <= X"5AC4C663";
    when 16#116A# => romdata <= X"12E8B79F";
    when 16#116B# => romdata <= X"0B92279A";
    when 16#116C# => romdata <= X"C7EF1936";
    when 16#116D# => romdata <= X"BCC30802";
    when 16#116E# => romdata <= X"B83DB3D1";
    when 16#116F# => romdata <= X"13BEF644";
    when 16#1170# => romdata <= X"52CAD7AC";
    when 16#1171# => romdata <= X"F6674FDA";
    when 16#1172# => romdata <= X"44023A66";
    when 16#1173# => romdata <= X"1019841A";
    when 16#1174# => romdata <= X"101BE80F";
    when 16#1175# => romdata <= X"DA4E3210";
    when 16#1176# => romdata <= X"AE774E43";
    when 16#1177# => romdata <= X"3A9ABD97";
    when 16#1178# => romdata <= X"F2755259";
    when 16#1179# => romdata <= X"AECE21F7";
    when 16#117A# => romdata <= X"A8C3B1A3";
    when 16#117B# => romdata <= X"D471F874";
    when 16#117C# => romdata <= X"D2EEC85B";
    when 16#117D# => romdata <= X"9B21BC0C";
    when 16#117E# => romdata <= X"2E2EC901";
    when 16#117F# => romdata <= X"6F847C60";
    when 16#1180# => romdata <= X"EE38BAF6";
    when 16#1181# => romdata <= X"F61704B0";
    when 16#1182# => romdata <= X"1509B521";
    when 16#1183# => romdata <= X"0A0534E4";
    when 16#1184# => romdata <= X"702F9319";
    when 16#1185# => romdata <= X"0C392E74";
    when 16#1186# => romdata <= X"9869B557";
    when 16#1187# => romdata <= X"2BB7AC4D";
    when 16#1188# => romdata <= X"7120E2BE";
    when 16#1189# => romdata <= X"CD6618CD";
    when 16#118A# => romdata <= X"376C4C1B";
    when 16#118B# => romdata <= X"4965F7D9";
    when 16#118C# => romdata <= X"D7340082";
    when 16#118D# => romdata <= X"4E88A5C7";
    when 16#118E# => romdata <= X"B5B66BA8";
    when 16#118F# => romdata <= X"8C3E0065";
    when 16#1190# => romdata <= X"F9628A9A";
    when 16#1191# => romdata <= X"C6B91A18";
    when 16#1192# => romdata <= X"82192FC5";
    when 16#1193# => romdata <= X"53E31403";
    when 16#1194# => romdata <= X"49934D20";
    when 16#1195# => romdata <= X"698C9F29";
    when 16#1196# => romdata <= X"1B537094";
    when 16#1197# => romdata <= X"8AF6CC90";
    when 16#1198# => romdata <= X"C837B9F3";
    when 16#1199# => romdata <= X"607F13CA";
    when 16#119A# => romdata <= X"FD492CEF";
    when 16#119B# => romdata <= X"1723376E";
    when 16#119C# => romdata <= X"6A5B813A";
    when 16#119D# => romdata <= X"56301B88";
    when 16#119E# => romdata <= X"A8799519";
    when 16#119F# => romdata <= X"CB7646F3";
    when 16#11A0# => romdata <= X"3F91C44C";
    when 16#11A1# => romdata <= X"DBE7F768";
    when 16#11A2# => romdata <= X"D7DD9B32";
    when 16#11A3# => romdata <= X"3A5002D2";
    when 16#11A4# => romdata <= X"F784C410";
    when 16#11A5# => romdata <= X"1AF90D6E";
    when 16#11A6# => romdata <= X"4C5ADE7D";
    when 16#11A7# => romdata <= X"085C79E8";
    when 16#11A8# => romdata <= X"27D43E10";
    when 16#11A9# => romdata <= X"DF63AC70";
    when 16#11AA# => romdata <= X"BCDF13DC";
    when 16#11AB# => romdata <= X"E0471B48";
    when 16#11AC# => romdata <= X"7C5ECB75";
    when 16#11AD# => romdata <= X"2B9C3E20";
    when 16#11AE# => romdata <= X"F75DBD24";
    when 16#11AF# => romdata <= X"3790C913";
    when 16#11B0# => romdata <= X"55ADFD71";
    when 16#11B1# => romdata <= X"99081BFE";
    when 16#11B2# => romdata <= X"A03D80E8";
    when 16#11B3# => romdata <= X"2445EC28";
    when 16#11B4# => romdata <= X"31FB5014";
    when 16#11B5# => romdata <= X"B85EFC2A";
    when 16#11B6# => romdata <= X"52748A8A";
    when 16#11B7# => romdata <= X"BFAC1BA3";
    when 16#11B8# => romdata <= X"904E178D";
    when 16#11B9# => romdata <= X"FBAB26C1";
    when 16#11BA# => romdata <= X"750228C9";
    when 16#11BB# => romdata <= X"A031104F";
    when 16#11BC# => romdata <= X"58BB3B91";
    when 16#11BD# => romdata <= X"905EDB9E";
    when 16#11BE# => romdata <= X"ADF7B0F6";
    when 16#11BF# => romdata <= X"DF22ACEB";
    when 16#11C0# => romdata <= X"0DE944E2";
    when 16#11C1# => romdata <= X"77809D77";
    when 16#11C2# => romdata <= X"507D18EA";
    when 16#11C3# => romdata <= X"EDAA1767";
    when 16#11C4# => romdata <= X"69739842";
    when 16#11C5# => romdata <= X"1115D04A";
    when 16#11C6# => romdata <= X"B2EBFC46";
    when 16#11C7# => romdata <= X"6E99F0AA";
    when 16#11C8# => romdata <= X"540482A4";
    when 16#11C9# => romdata <= X"9C6AC8FF";
    when 16#11CA# => romdata <= X"95E3F962";
    when 16#11CB# => romdata <= X"734B03EF";
    when 16#11CC# => romdata <= X"39873A93";
    when 16#11CD# => romdata <= X"B70470B4";
    when 16#11CE# => romdata <= X"6FFFDFDC";
    when 16#11CF# => romdata <= X"15C89F8F";
    when 16#11D0# => romdata <= X"E2F4637B";
    when 16#11D1# => romdata <= X"59F9BF9C";
    when 16#11D2# => romdata <= X"5752D9F8";
    when 16#11D3# => romdata <= X"AE7EA75D";
    when 16#11D4# => romdata <= X"1EAF1C22";
    when 16#11D5# => romdata <= X"CA27E5D5";
    when 16#11D6# => romdata <= X"C9499624";
    when 16#11D7# => romdata <= X"105D61BE";
    when 16#11D8# => romdata <= X"2A691F91";
    when 16#11D9# => romdata <= X"94D27741";
    when 16#11DA# => romdata <= X"4532A5E6";
    when 16#11DB# => romdata <= X"C63875F7";
    when 16#11DC# => romdata <= X"F20DD13C";
    when 16#11DD# => romdata <= X"6EE73B0C";
    when 16#11DE# => romdata <= X"3568392B";
    when 16#11DF# => romdata <= X"14A50428";
    when 16#11E0# => romdata <= X"43926472";
    when 16#11E1# => romdata <= X"ABA343D2";
    when 16#11E2# => romdata <= X"C4277921";
    when 16#11E3# => romdata <= X"99B543BE";
    when 16#11E4# => romdata <= X"1D43A178";
    when 16#11E5# => romdata <= X"FAA7ECF5";
    when 16#11E6# => romdata <= X"3B98AB75";
    when 16#11E7# => romdata <= X"28D8E1B8";
    when 16#11E8# => romdata <= X"B82C52D9";
    when 16#11E9# => romdata <= X"73CA0427";
    when 16#11EA# => romdata <= X"63650583";
    when 16#11EB# => romdata <= X"7F94284E";
    when 16#11EC# => romdata <= X"8D6B4F49";
    when 16#11ED# => romdata <= X"6FC5A48B";
    when 16#11EE# => romdata <= X"7958D468";
    when 16#11EF# => romdata <= X"1DA00651";
    when 16#11F0# => romdata <= X"B8A7BC56";
    when 16#11F1# => romdata <= X"EC859C07";
    when 16#11F2# => romdata <= X"1E4396A0";
    when 16#11F3# => romdata <= X"5F33588B";
    when 16#11F4# => romdata <= X"8087EFE9";
    when 16#11F5# => romdata <= X"635E565E";
    when 16#11F6# => romdata <= X"6B5A8A70";
    when 16#11F7# => romdata <= X"DA70F50E";
    when 16#11F8# => romdata <= X"CAD1A85E";
    when 16#11F9# => romdata <= X"6E36FF07";
    when 16#11FA# => romdata <= X"B4FB3B91";
    when 16#11FB# => romdata <= X"19EDE0B6";
    when 16#11FC# => romdata <= X"11CFA91D";
    when 16#11FD# => romdata <= X"9D4C58C1";
    when 16#11FE# => romdata <= X"F4815B07";
    when 16#11FF# => romdata <= X"B9EB1DE0";
    when 16#1200# => romdata <= X"CD37D0FB";
    when 16#1201# => romdata <= X"0043D034";
    when 16#1202# => romdata <= X"44A939E9";
    when 16#1203# => romdata <= X"3676B9DA";
    when 16#1204# => romdata <= X"F5F2D19A";
    when 16#1205# => romdata <= X"2615E3D9";
    when 16#1206# => romdata <= X"7D624E62";
    when 16#1207# => romdata <= X"ACAC8098";
    when 16#1208# => romdata <= X"099FDB9A";
    when 16#1209# => romdata <= X"5A2F4B3A";
    when 16#120A# => romdata <= X"CF20F75B";
    when 16#120B# => romdata <= X"6807A5A3";
    when 16#120C# => romdata <= X"F157C2C0";
    when 16#120D# => romdata <= X"F479158F";
    when 16#120E# => romdata <= X"4A10FB49";
    when 16#120F# => romdata <= X"72855F3A";
    when 16#1210# => romdata <= X"E2FDCBDE";
    when 16#1211# => romdata <= X"EC00A4D4";
    when 16#1212# => romdata <= X"70AADF5F";
    when 16#1213# => romdata <= X"5E571818";
    when 16#1214# => romdata <= X"AD6E872D";
    when 16#1215# => romdata <= X"897E2DDC";
    when 16#1216# => romdata <= X"40200696";
    when 16#1217# => romdata <= X"5ADF1658";
    when 16#1218# => romdata <= X"2B1E06B1";
    when 16#1219# => romdata <= X"861BF7D0";
    when 16#121A# => romdata <= X"C7E7BA49";
    when 16#121B# => romdata <= X"1C79E862";
    when 16#121C# => romdata <= X"24AF6B24";
    when 16#121D# => romdata <= X"6317F725";
    when 16#121E# => romdata <= X"FA74DD83";
    when 16#121F# => romdata <= X"76D63D79";
    when 16#1220# => romdata <= X"93FE2F2B";
    when 16#1221# => romdata <= X"BBB2F1DA";
    when 16#1222# => romdata <= X"9238C6F3";
    when 16#1223# => romdata <= X"FFCAEC50";
    when 16#1224# => romdata <= X"FF61E645";
    when 16#1225# => romdata <= X"FADEB6E0";
    when 16#1226# => romdata <= X"3F883892";
    when 16#1227# => romdata <= X"C42CCCF9";
    when 16#1228# => romdata <= X"04708B12";
    when 16#1229# => romdata <= X"3C9271A6";
    when 16#122A# => romdata <= X"70D4DCFC";
    when 16#122B# => romdata <= X"D602951D";
    when 16#122C# => romdata <= X"12F52139";
    when 16#122D# => romdata <= X"37CA2C05";
    when 16#122E# => romdata <= X"ADDE9EE3";
    when 16#122F# => romdata <= X"908E99AA";
    when 16#1230# => romdata <= X"E8DA3195";
    when 16#1231# => romdata <= X"1C36D36D";
    when 16#1232# => romdata <= X"671CD7BF";
    when 16#1233# => romdata <= X"15DF60B7";
    when 16#1234# => romdata <= X"07F00BF6";
    when 16#1235# => romdata <= X"EBBE5476";
    when 16#1236# => romdata <= X"926D0156";
    when 16#1237# => romdata <= X"28A85758";
    when 16#1238# => romdata <= X"BFF35C4A";
    when 16#1239# => romdata <= X"C540F39E";
    when 16#123A# => romdata <= X"761B2ED3";
    when 16#123B# => romdata <= X"CA9116E8";
    when 16#123C# => romdata <= X"680E28BC";
    when 16#123D# => romdata <= X"387058E0";
    when 16#123E# => romdata <= X"F69345CC";
    when 16#123F# => romdata <= X"6AB3AD16";
    when 16#1240# => romdata <= X"0E9F2BC4";
    when 16#1241# => romdata <= X"D6047A19";
    when 16#1242# => romdata <= X"34E15D3D";
    when 16#1243# => romdata <= X"7A242A29";
    when 16#1244# => romdata <= X"6333C092";
    when 16#1245# => romdata <= X"96981BBF";
    when 16#1246# => romdata <= X"3B8577E4";
    when 16#1247# => romdata <= X"B8ED2A36";
    when 16#1248# => romdata <= X"24866111";
    when 16#1249# => romdata <= X"F6638F89";
    when 16#124A# => romdata <= X"55431195";
    when 16#124B# => romdata <= X"B60C5C08";
    when 16#124C# => romdata <= X"9F9897DD";
    when 16#124D# => romdata <= X"F0D34A3D";
    when 16#124E# => romdata <= X"C627CE33";
    when 16#124F# => romdata <= X"7AC8128C";
    when 16#1250# => romdata <= X"28B63A39";
    when 16#1251# => romdata <= X"4908E4C0";
    when 16#1252# => romdata <= X"83BCC452";
    when 16#1253# => romdata <= X"2DB8CE57";
    when 16#1254# => romdata <= X"20C45EF7";
    when 16#1255# => romdata <= X"6B271622";
    when 16#1256# => romdata <= X"5E53405F";
    when 16#1257# => romdata <= X"CAAAA72A";
    when 16#1258# => romdata <= X"C1982265";
    when 16#1259# => romdata <= X"75D52251";
    when 16#125A# => romdata <= X"95F106C1";
    when 16#125B# => romdata <= X"249E4B87";
    when 16#125C# => romdata <= X"AC05287A";
    when 16#125D# => romdata <= X"3ABE6C51";
    when 16#125E# => romdata <= X"A2A41E07";
    when 16#125F# => romdata <= X"F56ECDC4";
    when 16#1260# => romdata <= X"6E989A85";
    when 16#1261# => romdata <= X"68D35669";
    when 16#1262# => romdata <= X"B525A6FF";
    when 16#1263# => romdata <= X"CA90DC91";
    when 16#1264# => romdata <= X"D3013967";
    when 16#1265# => romdata <= X"F6A5F4C0";
    when 16#1266# => romdata <= X"22FFCC17";
    when 16#1267# => romdata <= X"751B68FB";
    when 16#1268# => romdata <= X"0D8F16FC";
    when 16#1269# => romdata <= X"9229851D";
    when 16#126A# => romdata <= X"FDCC0608";
    when 16#126B# => romdata <= X"38F923BD";
    when 16#126C# => romdata <= X"44C1AD70";
    when 16#126D# => romdata <= X"A993E8EB";
    when 16#126E# => romdata <= X"AC1667DA";
    when 16#126F# => romdata <= X"80F91B66";
    when 16#1270# => romdata <= X"F8F5B375";
    when 16#1271# => romdata <= X"D3527518";
    when 16#1272# => romdata <= X"8E3C7702";
    when 16#1273# => romdata <= X"C2312CEA";
    when 16#1274# => romdata <= X"C5B20D67";
    when 16#1275# => romdata <= X"BB344004";
    when 16#1276# => romdata <= X"01BDF1DB";
    when 16#1277# => romdata <= X"FE79DFA0";
    when 16#1278# => romdata <= X"EB73F173";
    when 16#1279# => romdata <= X"A0480721";
    when 16#127A# => romdata <= X"5DA5CE8E";
    when 16#127B# => romdata <= X"1D28F212";
    when 16#127C# => romdata <= X"6424C3DB";
    when 16#127D# => romdata <= X"44ADCD7A";
    when 16#127E# => romdata <= X"961260FD";
    when 16#127F# => romdata <= X"BCAB31E0";
    when 16#1280# => romdata <= X"CAA02DD1";
    when 16#1281# => romdata <= X"9DB9C721";
    when 16#1282# => romdata <= X"EB35AB7D";
    when 16#1283# => romdata <= X"64B8A387";
    when 16#1284# => romdata <= X"79642724";
    when 16#1285# => romdata <= X"2698A47D";
    when 16#1286# => romdata <= X"832C3F1A";
    when 16#1287# => romdata <= X"D4DDA0B5";
    when 16#1288# => romdata <= X"926FFCE9";
    when 16#1289# => romdata <= X"319EEEDA";
    when 16#128A# => romdata <= X"1565ECB0";
    when 16#128B# => romdata <= X"FA1EEDB4";
    when 16#128C# => romdata <= X"24414120";
    when 16#128D# => romdata <= X"AAE8CFD0";
    when 16#128E# => romdata <= X"BE88D4D2";
    when 16#128F# => romdata <= X"48899A0B";
    when 16#1290# => romdata <= X"CE31F9BE";
    when 16#1291# => romdata <= X"E7A4DC4D";
    when 16#1292# => romdata <= X"B3C3B104";
    when 16#1293# => romdata <= X"44FAD6AD";
    when 16#1294# => romdata <= X"CCE28F0E";
    when 16#1295# => romdata <= X"DF7B8085";
    when 16#1296# => romdata <= X"36ACF5EB";
    when 16#1297# => romdata <= X"05AADAE9";
    when 16#1298# => romdata <= X"2693EE02";
    when 16#1299# => romdata <= X"C9512B3E";
    when 16#129A# => romdata <= X"EF000844";
    when 16#129B# => romdata <= X"BA35E246";
    when 16#129C# => romdata <= X"20A2E893";
    when 16#129D# => romdata <= X"5354B843";
    when 16#129E# => romdata <= X"2C07C8FD";
    when 16#129F# => romdata <= X"615534BC";
    when 16#12A0# => romdata <= X"FD0D8E3B";
    when 16#12A1# => romdata <= X"572BF2CF";
    when 16#12A2# => romdata <= X"06AD3439";
    when 16#12A3# => romdata <= X"97590FE8";
    when 16#12A4# => romdata <= X"B244A32B";
    when 16#12A5# => romdata <= X"BE69125B";
    when 16#12A6# => romdata <= X"5D7C5E51";
    when 16#12A7# => romdata <= X"3A493724";
    when 16#12A8# => romdata <= X"EEA8DA6C";
    when 16#12A9# => romdata <= X"B0FFF3AC";
    when 16#12AA# => romdata <= X"F1C5085A";
    when 16#12AB# => romdata <= X"8120694C";
    when 16#12AC# => romdata <= X"BC40FAE1";
    when 16#12AD# => romdata <= X"A6326FD7";
    when 16#12AE# => romdata <= X"1487CC3B";
    when 16#12AF# => romdata <= X"E7C10A34";
    when 16#12B0# => romdata <= X"315CDFFA";
    when 16#12B1# => romdata <= X"8C618B68";
    when 16#12B2# => romdata <= X"EA93D330";
    when 16#12B3# => romdata <= X"945586B0";
    when 16#12B4# => romdata <= X"80381F00";
    when 16#12B5# => romdata <= X"76351B88";
    when 16#12B6# => romdata <= X"8087F56B";
    when 16#12B7# => romdata <= X"969E6D6A";
    when 16#12B8# => romdata <= X"311AE03C";
    when 16#12B9# => romdata <= X"C79FF686";
    when 16#12BA# => romdata <= X"1E715C9D";
    when 16#12BB# => romdata <= X"A9AEE751";
    when 16#12BC# => romdata <= X"F1220661";
    when 16#12BD# => romdata <= X"581C75DC";
    when 16#12BE# => romdata <= X"EC0515A1";
    when 16#12BF# => romdata <= X"C9259B9C";
    when 16#12C0# => romdata <= X"F8E944CE";
    when 16#12C1# => romdata <= X"C4B1754E";
    when 16#12C2# => romdata <= X"5809E985";
    when 16#12C3# => romdata <= X"D6F43FE4";
    when 16#12C4# => romdata <= X"57108932";
    when 16#12C5# => romdata <= X"42ADE0D3";
    when 16#12C6# => romdata <= X"B84F1E19";
    when 16#12C7# => romdata <= X"42B7A956";
    when 16#12C8# => romdata <= X"48611595";
    when 16#12C9# => romdata <= X"FED13F54";
    when 16#12CA# => romdata <= X"6CA11DB8";
    when 16#12CB# => romdata <= X"E5A55A3C";
    when 16#12CC# => romdata <= X"3C78C379";
    when 16#12CD# => romdata <= X"3C6689E1";
    when 16#12CE# => romdata <= X"B3AFB5F6";
    when 16#12CF# => romdata <= X"7526A480";
    when 16#12D0# => romdata <= X"DF923A58";
    when 16#12D1# => romdata <= X"6A779F94";
    when 16#12D2# => romdata <= X"A09CF963";
    when 16#12D3# => romdata <= X"594FF4B0";
    when 16#12D4# => romdata <= X"A387876E";
    when 16#12D5# => romdata <= X"BB3E8FAB";
    when 16#12D6# => romdata <= X"888C97F6";
    when 16#12D7# => romdata <= X"773E7F03";
    when 16#12D8# => romdata <= X"17B038E4";
    when 16#12D9# => romdata <= X"7DD7D109";
    when 16#12DA# => romdata <= X"545BB072";
    when 16#12DB# => romdata <= X"63B1AA84";
    when 16#12DC# => romdata <= X"284B86E4";
    when 16#12DD# => romdata <= X"7FFB9784";
    when 16#12DE# => romdata <= X"A171D101";
    when 16#12DF# => romdata <= X"E7B0A6D3";
    when 16#12E0# => romdata <= X"8BCAE7E6";
    when 16#12E1# => romdata <= X"3D827C99";
    when 16#12E2# => romdata <= X"9BF55172";
    when 16#12E3# => romdata <= X"8FFC642E";
    when 16#12E4# => romdata <= X"E690B01D";
    when 16#12E5# => romdata <= X"486CB6EB";
    when 16#12E6# => romdata <= X"EEB9D5C8";
    when 16#12E7# => romdata <= X"88112589";
    when 16#12E8# => romdata <= X"EA5CBC9B";
    when 16#12E9# => romdata <= X"DF49E675";
    when 16#12EA# => romdata <= X"96522341";
    when 16#12EB# => romdata <= X"6D6DA02D";
    when 16#12EC# => romdata <= X"2333BFD4";
    when 16#12ED# => romdata <= X"614706BF";
    when 16#12EE# => romdata <= X"13373973";
    when 16#12EF# => romdata <= X"207C849A";
    when 16#12F0# => romdata <= X"0DE41EBA";
    when 16#12F1# => romdata <= X"137FDF79";
    when 16#12F2# => romdata <= X"A1EB25D7";
    when 16#12F3# => romdata <= X"4E30CF60";
    when 16#12F4# => romdata <= X"B577C278";
    when 16#12F5# => romdata <= X"7DF04740";
    when 16#12F6# => romdata <= X"BA8CADE3";
    when 16#12F7# => romdata <= X"F9DA55D3";
    when 16#12F8# => romdata <= X"F0084F02";
    when 16#12F9# => romdata <= X"809E3754";
    when 16#12FA# => romdata <= X"3239E0A7";
    when 16#12FB# => romdata <= X"1E99751E";
    when 16#12FC# => romdata <= X"EB21CB3B";
    when 16#12FD# => romdata <= X"41488244";
    when 16#12FE# => romdata <= X"193A4868";
    when 16#12FF# => romdata <= X"CBA92760";
    when 16#1300# => romdata <= X"FB227530";
    when 16#1301# => romdata <= X"F82BD527";
    when 16#1302# => romdata <= X"E648619E";
    when 16#1303# => romdata <= X"532D7646";
    when 16#1304# => romdata <= X"A5ABBD15";
    when 16#1305# => romdata <= X"DB91A6E7";
    when 16#1306# => romdata <= X"033DFECC";
    when 16#1307# => romdata <= X"C65D095A";
    when 16#1308# => romdata <= X"3D83AB77";
    when 16#1309# => romdata <= X"EDD2F3FE";
    when 16#130A# => romdata <= X"C52659CB";
    when 16#130B# => romdata <= X"3AD1BEB0";
    when 16#130C# => romdata <= X"09D7A1C9";
    when 16#130D# => romdata <= X"BFB54429";
    when 16#130E# => romdata <= X"1EC1C67B";
    when 16#130F# => romdata <= X"75DD6DAB";
    when 16#1310# => romdata <= X"06E70C32";
    when 16#1311# => romdata <= X"C7149831";
    when 16#1312# => romdata <= X"39DE4A41";
    when 16#1313# => romdata <= X"EE07B4F3";
    when 16#1314# => romdata <= X"C03BF566";
    when 16#1315# => romdata <= X"558484F1";
    when 16#1316# => romdata <= X"9A3BB674";
    when 16#1317# => romdata <= X"B6795F0D";
    when 16#1318# => romdata <= X"8537BC31";
    when 16#1319# => romdata <= X"BC8D7A38";
    when 16#131A# => romdata <= X"B2FF1B2E";
    when 16#131B# => romdata <= X"C8B78539";
    when 16#131C# => romdata <= X"B2251D0E";
    when 16#131D# => romdata <= X"385DE484";
    when 16#131E# => romdata <= X"B05A4114";
    when 16#131F# => romdata <= X"77681A3A";
    when 16#1320# => romdata <= X"E7527AC9";
    when 16#1321# => romdata <= X"8BC2943A";
    when 16#1322# => romdata <= X"F1CF7F09";
    when 16#1323# => romdata <= X"ACF2DDE4";
    when 16#1324# => romdata <= X"530AE896";
    when 16#1325# => romdata <= X"BDE1266F";
    when 16#1326# => romdata <= X"E916E833";
    when 16#1327# => romdata <= X"A1C0CAA2";
    when 16#1328# => romdata <= X"B2D2F598";
    when 16#1329# => romdata <= X"5AD47B2D";
    when 16#132A# => romdata <= X"0D1D3AFB";
    when 16#132B# => romdata <= X"6E50D4B3";
    when 16#132C# => romdata <= X"DA7DEEC4";
    when 16#132D# => romdata <= X"385E6CA8";
    when 16#132E# => romdata <= X"FE22760F";
    when 16#132F# => romdata <= X"92807AC5";
    when 16#1330# => romdata <= X"5556AAF7";
    when 16#1331# => romdata <= X"973E8016";
    when 16#1332# => romdata <= X"ADFD43A3";
    when 16#1333# => romdata <= X"919088B7";
    when 16#1334# => romdata <= X"68351B10";
    when 16#1335# => romdata <= X"57498D2D";
    when 16#1336# => romdata <= X"668D7C1E";
    when 16#1337# => romdata <= X"8C634380";
    when 16#1338# => romdata <= X"55FDF7D3";
    when 16#1339# => romdata <= X"6C5E7DF0";
    when 16#133A# => romdata <= X"2FCAFCBD";
    when 16#133B# => romdata <= X"9291A214";
    when 16#133C# => romdata <= X"9E7B429B";
    when 16#133D# => romdata <= X"3202D329";
    when 16#133E# => romdata <= X"E47CED51";
    when 16#133F# => romdata <= X"EA577177";
    when 16#1340# => romdata <= X"2E308C5B";
    when 16#1341# => romdata <= X"EBA7B934";
    when 16#1342# => romdata <= X"597540D8";
    when 16#1343# => romdata <= X"3DBEC6C3";
    when 16#1344# => romdata <= X"BC61A96E";
    when 16#1345# => romdata <= X"A4CB2D75";
    when 16#1346# => romdata <= X"30D9D760";
    when 16#1347# => romdata <= X"AA940333";
    when 16#1348# => romdata <= X"8CD95B82";
    when 16#1349# => romdata <= X"9F17547C";
    when 16#134A# => romdata <= X"5A90D161";
    when 16#134B# => romdata <= X"F7B8CE00";
    when 16#134C# => romdata <= X"37EBF403";
    when 16#134D# => romdata <= X"C91C0D0C";
    when 16#134E# => romdata <= X"70C589BA";
    when 16#134F# => romdata <= X"87CAE8DF";
    when 16#1350# => romdata <= X"26CF1428";
    when 16#1351# => romdata <= X"1E235A68";
    when 16#1352# => romdata <= X"6CCD10E2";
    when 16#1353# => romdata <= X"D520A762";
    when 16#1354# => romdata <= X"65C4C278";
    when 16#1355# => romdata <= X"0EDFD070";
    when 16#1356# => romdata <= X"5E89EFE3";
    when 16#1357# => romdata <= X"C953FE76";
    when 16#1358# => romdata <= X"0DE45A8C";
    when 16#1359# => romdata <= X"F1F2D3F3";
    when 16#135A# => romdata <= X"6DE3164D";
    when 16#135B# => romdata <= X"5BC2CF32";
    when 16#135C# => romdata <= X"204228AD";
    when 16#135D# => romdata <= X"D7C182EC";
    when 16#135E# => romdata <= X"55F1158A";
    when 16#135F# => romdata <= X"FA9358BE";
    when 16#1360# => romdata <= X"179C722A";
    when 16#1361# => romdata <= X"DAF1D0BF";
    when 16#1362# => romdata <= X"1306A0B5";
    when 16#1363# => romdata <= X"6218857F";
    when 16#1364# => romdata <= X"C5C21001";
    when 16#1365# => romdata <= X"499F61E2";
    when 16#1366# => romdata <= X"73442281";
    when 16#1367# => romdata <= X"E585B3E6";
    when 16#1368# => romdata <= X"DCE148AA";
    when 16#1369# => romdata <= X"97B6622B";
    when 16#136A# => romdata <= X"23BDAECF";
    when 16#136B# => romdata <= X"983BF186";
    when 16#136C# => romdata <= X"F1B34962";
    when 16#136D# => romdata <= X"764758AC";
    when 16#136E# => romdata <= X"3C20C840";
    when 16#136F# => romdata <= X"36061D49";
    when 16#1370# => romdata <= X"CA33B3C3";
    when 16#1371# => romdata <= X"FCDF03F4";
    when 16#1372# => romdata <= X"7F7E53B9";
    when 16#1373# => romdata <= X"40DBB6E1";
    when 16#1374# => romdata <= X"E4A26702";
    when 16#1375# => romdata <= X"A118E525";
    when 16#1376# => romdata <= X"A9A0EC22";
    when 16#1377# => romdata <= X"9085C925";
    when 16#1378# => romdata <= X"D133750E";
    when 16#1379# => romdata <= X"D0B200CB";
    when 16#137A# => romdata <= X"28A11328";
    when 16#137B# => romdata <= X"9DE143D1";
    when 16#137C# => romdata <= X"D5839D2A";
    when 16#137D# => romdata <= X"F8B0525E";
    when 16#137E# => romdata <= X"0027F34F";
    when 16#137F# => romdata <= X"F32106A0";
    when 16#1380# => romdata <= X"9E5DA18A";
    when 16#1381# => romdata <= X"19514CCC";
    when 16#1382# => romdata <= X"849E9697";
    when 16#1383# => romdata <= X"AE4BD1B3";
    when 16#1384# => romdata <= X"17BB3492";
    when 16#1385# => romdata <= X"7D0461A9";
    when 16#1386# => romdata <= X"6A7AF4A5";
    when 16#1387# => romdata <= X"D6C13107";
    when 16#1388# => romdata <= X"FFB9DE38";
    when 16#1389# => romdata <= X"C5E8CB7C";
    when 16#138A# => romdata <= X"5682827F";
    when 16#138B# => romdata <= X"57D94ED2";
    when 16#138C# => romdata <= X"E77D36F9";
    when 16#138D# => romdata <= X"F1CB05E4";
    when 16#138E# => romdata <= X"C2C62B1D";
    when 16#138F# => romdata <= X"E254C7B1";
    when 16#1390# => romdata <= X"CB236FC4";
    when 16#1391# => romdata <= X"ED70BF8D";
    when 16#1392# => romdata <= X"D1F43AC7";
    when 16#1393# => romdata <= X"73C16A37";
    when 16#1394# => romdata <= X"392B895F";
    when 16#1395# => romdata <= X"8B157578";
    when 16#1396# => romdata <= X"C477C85E";
    when 16#1397# => romdata <= X"53FA7CA5";
    when 16#1398# => romdata <= X"8BE70D91";
    when 16#1399# => romdata <= X"87AF5F7A";
    when 16#139A# => romdata <= X"18D5A1E5";
    when 16#139B# => romdata <= X"642335E4";
    when 16#139C# => romdata <= X"6C2F8F46";
    when 16#139D# => romdata <= X"91AEEE6A";
    when 16#139E# => romdata <= X"9692E21B";
    when 16#139F# => romdata <= X"9668E2C0";
    when 16#13A0# => romdata <= X"83D9F45C";
    when 16#13A1# => romdata <= X"2DB3E991";
    when 16#13A2# => romdata <= X"588BA87A";
    when 16#13A3# => romdata <= X"0A238087";
    when 16#13A4# => romdata <= X"32EE39E8";
    when 16#13A5# => romdata <= X"B3C876BE";
    when 16#13A6# => romdata <= X"79227C78";
    when 16#13A7# => romdata <= X"2F07EE3F";
    when 16#13A8# => romdata <= X"B3086AF9";
    when 16#13A9# => romdata <= X"13D71D71";
    when 16#13AA# => romdata <= X"910A0F56";
    when 16#13AB# => romdata <= X"D62B5DE5";
    when 16#13AC# => romdata <= X"E224F785";
    when 16#13AD# => romdata <= X"6A42A4A1";
    when 16#13AE# => romdata <= X"B2AFE380";
    when 16#13AF# => romdata <= X"827BE86E";
    when 16#13B0# => romdata <= X"381FCE48";
    when 16#13B1# => romdata <= X"6FD08A91";
    when 16#13B2# => romdata <= X"B22BD91D";
    when 16#13B3# => romdata <= X"09615F41";
    when 16#13B4# => romdata <= X"7E178C55";
    when 16#13B5# => romdata <= X"93E41B09";
    when 16#13B6# => romdata <= X"17E07513";
    when 16#13B7# => romdata <= X"3960AD28";
    when 16#13B8# => romdata <= X"B4DD4096";
    when 16#13B9# => romdata <= X"D1E84BEF";
    when 16#13BA# => romdata <= X"1363098D";
    when 16#13BB# => romdata <= X"DE92C29C";
    when 16#13BC# => romdata <= X"D508C40B";
    when 16#13BD# => romdata <= X"A7E785F4";
    when 16#13BE# => romdata <= X"6C1E0DC7";
    when 16#13BF# => romdata <= X"2E729D39";
    when 16#13C0# => romdata <= X"4911DA91";
    when 16#13C1# => romdata <= X"9EA6F94D";
    when 16#13C2# => romdata <= X"14567FFA";
    when 16#13C3# => romdata <= X"DC61CEB8";
    when 16#13C4# => romdata <= X"DCA2821B";
    when 16#13C5# => romdata <= X"1CF04847";
    when 16#13C6# => romdata <= X"7E2433E9";
    when 16#13C7# => romdata <= X"DC718DE6";
    when 16#13C8# => romdata <= X"18EDEEF3";
    when 16#13C9# => romdata <= X"02CDCB5D";
    when 16#13CA# => romdata <= X"E472656D";
    when 16#13CB# => romdata <= X"6687DC41";
    when 16#13CC# => romdata <= X"EA34C2BB";
    when 16#13CD# => romdata <= X"4DF1CA08";
    when 16#13CE# => romdata <= X"DCB933BE";
    when 16#13CF# => romdata <= X"3EF4B419";
    when 16#13D0# => romdata <= X"158BA0B6";
    when 16#13D1# => romdata <= X"8AE82A64";
    when 16#13D2# => romdata <= X"ADD58559";
    when 16#13D3# => romdata <= X"214FD88A";
    when 16#13D4# => romdata <= X"4CB34D99";
    when 16#13D5# => romdata <= X"F6463106";
    when 16#13D6# => romdata <= X"97DA982C";
    when 16#13D7# => romdata <= X"2FD4EE06";
    when 16#13D8# => romdata <= X"9DC1CB10";
    when 16#13D9# => romdata <= X"2125C34A";
    when 16#13DA# => romdata <= X"89AB20F1";
    when 16#13DB# => romdata <= X"7B6EF648";
    when 16#13DC# => romdata <= X"A8346273";
    when 16#13DD# => romdata <= X"20410FF6";
    when 16#13DE# => romdata <= X"881C7919";
    when 16#13DF# => romdata <= X"AE4E71CB";
    when 16#13E0# => romdata <= X"AE5F8200";
    when 16#13E1# => romdata <= X"E523934D";
    when 16#13E2# => romdata <= X"84BFA897";
    when 16#13E3# => romdata <= X"C44B89B9";
    when 16#13E4# => romdata <= X"BC6BC012";
    when 16#13E5# => romdata <= X"9F7F97EE";
    when 16#13E6# => romdata <= X"0EC049BA";
    when 16#13E7# => romdata <= X"1AFD67D0";
    when 16#13E8# => romdata <= X"0CD624A7";
    when 16#13E9# => romdata <= X"5FF5A305";
    when 16#13EA# => romdata <= X"14399BE4";
    when 16#13EB# => romdata <= X"801CED05";
    when 16#13EC# => romdata <= X"7B498B9D";
    when 16#13ED# => romdata <= X"BBF0EB99";
    when 16#13EE# => romdata <= X"44295D5B";
    when 16#13EF# => romdata <= X"6AE968C4";
    when 16#13F0# => romdata <= X"B8BBD2B9";
    when 16#13F1# => romdata <= X"A9E17A30";
    when 16#13F2# => romdata <= X"39C5FA35";
    when 16#13F3# => romdata <= X"A0D30AA5";
    when 16#13F4# => romdata <= X"4CA426C5";
    when 16#13F5# => romdata <= X"8353943D";
    when 16#13F6# => romdata <= X"DDD3FD18";
    when 16#13F7# => romdata <= X"5895C0DA";
    when 16#13F8# => romdata <= X"EE950455";
    when 16#13F9# => romdata <= X"FC131F52";
    when 16#13FA# => romdata <= X"0B46AE11";
    when 16#13FB# => romdata <= X"8C7406D0";
    when 16#13FC# => romdata <= X"A72BE612";
    when 16#13FD# => romdata <= X"7C530773";
    when 16#13FE# => romdata <= X"0AD441B6";
    when 16#13FF# => romdata <= X"FC3D1E00";
    when 16#1400# => romdata <= X"8589F839";
    when 16#1401# => romdata <= X"6F5B1C54";
    when 16#1402# => romdata <= X"CAF2B17D";
    when 16#1403# => romdata <= X"4C152CEF";
    when 16#1404# => romdata <= X"347E66EC";
    when 16#1405# => romdata <= X"7903C878";
    when 16#1406# => romdata <= X"F2823D4A";
    when 16#1407# => romdata <= X"DB9E7CCF";
    when 16#1408# => romdata <= X"AFEBB926";
    when 16#1409# => romdata <= X"B7EEB4AE";
    when 16#140A# => romdata <= X"1BECA339";
    when 16#140B# => romdata <= X"A027CE8E";
    when 16#140C# => romdata <= X"F9979575";
    when 16#140D# => romdata <= X"32FA871F";
    when 16#140E# => romdata <= X"356E0326";
    when 16#140F# => romdata <= X"ECE0BCE3";
    when 16#1410# => romdata <= X"399F8117";
    when 16#1411# => romdata <= X"9BF78C5C";
    when 16#1412# => romdata <= X"7D135018";
    when 16#1413# => romdata <= X"ABC340C0";
    when 16#1414# => romdata <= X"BE58D306";
    when 16#1415# => romdata <= X"3DD7CDA4";
    when 16#1416# => romdata <= X"C1918A01";
    when 16#1417# => romdata <= X"87BACF83";
    when 16#1418# => romdata <= X"0C8B6900";
    when 16#1419# => romdata <= X"D43B62E0";
    when 16#141A# => romdata <= X"4DF6E831";
    when 16#141B# => romdata <= X"CFEFA13B";
    when 16#141C# => romdata <= X"DB5E873A";
    when 16#141D# => romdata <= X"527F2432";
    when 16#141E# => romdata <= X"7C95DB4B";
    when 16#141F# => romdata <= X"BDB65C81";
    when 16#1420# => romdata <= X"A20F959F";
    when 16#1421# => romdata <= X"828F5DAE";
    when 16#1422# => romdata <= X"4DC13E5C";
    when 16#1423# => romdata <= X"AC7417EE";
    when 16#1424# => romdata <= X"089401FB";
    when 16#1425# => romdata <= X"497ABE10";
    when 16#1426# => romdata <= X"144E28EA";
    when 16#1427# => romdata <= X"383E61D4";
    when 16#1428# => romdata <= X"A9B63B61";
    when 16#1429# => romdata <= X"8AA7CEA4";
    when 16#142A# => romdata <= X"588B2911";
    when 16#142B# => romdata <= X"EC581F50";
    when 16#142C# => romdata <= X"6062B05E";
    when 16#142D# => romdata <= X"7BEF723A";
    when 16#142E# => romdata <= X"5A465C9F";
    when 16#142F# => romdata <= X"BE70E313";
    when 16#1430# => romdata <= X"753BDE31";
    when 16#1431# => romdata <= X"02845A79";
    when 16#1432# => romdata <= X"A206BF7D";
    when 16#1433# => romdata <= X"996F49A2";
    when 16#1434# => romdata <= X"1752D534";
    when 16#1435# => romdata <= X"B73EE83B";
    when 16#1436# => romdata <= X"48C1A225";
    when 16#1437# => romdata <= X"F85F5103";
    when 16#1438# => romdata <= X"DDB9B6B8";
    when 16#1439# => romdata <= X"380F61AA";
    when 16#143A# => romdata <= X"F26E5CA6";
    when 16#143B# => romdata <= X"43EB62EA";
    when 16#143C# => romdata <= X"F58AFEE0";
    when 16#143D# => romdata <= X"D3494E4F";
    when 16#143E# => romdata <= X"7A4F642A";
    when 16#143F# => romdata <= X"3454F4F5";
    when 16#1440# => romdata <= X"6A406A26";
    when 16#1441# => romdata <= X"4148FF5D";
    when 16#1442# => romdata <= X"AC9DF5F1";
    when 16#1443# => romdata <= X"51C12E89";
    when 16#1444# => romdata <= X"ED9D4FDC";
    when 16#1445# => romdata <= X"C04EC5F0";
    when 16#1446# => romdata <= X"022DF8CB";
    when 16#1447# => romdata <= X"AF3CBC67";
    when 16#1448# => romdata <= X"CED2853F";
    when 16#1449# => romdata <= X"B4F8C589";
    when 16#144A# => romdata <= X"4C96CD00";
    when 16#144B# => romdata <= X"550950E7";
    when 16#144C# => romdata <= X"EA2A26C8";
    when 16#144D# => romdata <= X"0A72DF53";
    when 16#144E# => romdata <= X"3270A0E2";
    when 16#144F# => romdata <= X"3EDBAA4D";
    when 16#1450# => romdata <= X"0BE935D6";
    when 16#1451# => romdata <= X"2CC885E1";
    when 16#1452# => romdata <= X"CCE653D6";
    when 16#1453# => romdata <= X"6C51E49C";
    when 16#1454# => romdata <= X"43952042";
    when 16#1455# => romdata <= X"E1B2D043";
    when 16#1456# => romdata <= X"BDA1CFFC";
    when 16#1457# => romdata <= X"1E98A3F8";
    when 16#1458# => romdata <= X"06EB587A";
    when 16#1459# => romdata <= X"4EC9AE29";
    when 16#145A# => romdata <= X"9BD838C6";
    when 16#145B# => romdata <= X"8B9BBF7C";
    when 16#145C# => romdata <= X"420C12B2";
    when 16#145D# => romdata <= X"3AA2793F";
    when 16#145E# => romdata <= X"A0248C93";
    when 16#145F# => romdata <= X"2A91BCDD";
    when 16#1460# => romdata <= X"641DCB38";
    when 16#1461# => romdata <= X"F0B2D718";
    when 16#1462# => romdata <= X"7D898692";
    when 16#1463# => romdata <= X"8DF4602B";
    when 16#1464# => romdata <= X"381BA13B";
    when 16#1465# => romdata <= X"26329113";
    when 16#1466# => romdata <= X"4628FC91";
    when 16#1467# => romdata <= X"C8EDE925";
    when 16#1468# => romdata <= X"94B39650";
    when 16#1469# => romdata <= X"B877D9A9";
    when 16#146A# => romdata <= X"1DAAA052";
    when 16#146B# => romdata <= X"95457DFB";
    when 16#146C# => romdata <= X"2C5D8207";
    when 16#146D# => romdata <= X"BBCDFE16";
    when 16#146E# => romdata <= X"AC5B9360";
    when 16#146F# => romdata <= X"0E33BC97";
    when 16#1470# => romdata <= X"0B38E188";
    when 16#1471# => romdata <= X"08B1A732";
    when 16#1472# => romdata <= X"88932035";
    when 16#1473# => romdata <= X"2B524B10";
    when 16#1474# => romdata <= X"9560136E";
    when 16#1475# => romdata <= X"605D3278";
    when 16#1476# => romdata <= X"4CA01F8B";
    when 16#1477# => romdata <= X"11D077C8";
    when 16#1478# => romdata <= X"1EAD6B7A";
    when 16#1479# => romdata <= X"5741C82D";
    when 16#147A# => romdata <= X"76CEEF76";
    when 16#147B# => romdata <= X"4FD07E36";
    when 16#147C# => romdata <= X"1D531B75";
    when 16#147D# => romdata <= X"106AF157";
    when 16#147E# => romdata <= X"2AD1375B";
    when 16#147F# => romdata <= X"2BBAB680";
    when 16#1480# => romdata <= X"A3E17A4C";
    when 16#1481# => romdata <= X"AD2ABE76";
    when 16#1482# => romdata <= X"E32D1850";
    when 16#1483# => romdata <= X"1899F8D6";
    when 16#1484# => romdata <= X"0D293BB1";
    when 16#1485# => romdata <= X"AC3ADB64";
    when 16#1486# => romdata <= X"F81148AF";
    when 16#1487# => romdata <= X"56741790";
    when 16#1488# => romdata <= X"F87F8B7A";
    when 16#1489# => romdata <= X"2D9A6E76";
    when 16#148A# => romdata <= X"45EA50B7";
    when 16#148B# => romdata <= X"5514C394";
    when 16#148C# => romdata <= X"508884CB";
    when 16#148D# => romdata <= X"F9E320B2";
    when 16#148E# => romdata <= X"4D41D824";
    when 16#148F# => romdata <= X"6EB3C163";
    when 16#1490# => romdata <= X"B9101240";
    when 16#1491# => romdata <= X"776C312D";
    when 16#1492# => romdata <= X"B63C3388";
    when 16#1493# => romdata <= X"9E3C1218";
    when 16#1494# => romdata <= X"43585047";
    when 16#1495# => romdata <= X"1C454486";
    when 16#1496# => romdata <= X"DF7FF4D2";
    when 16#1497# => romdata <= X"DC0AAA14";
    when 16#1498# => romdata <= X"980F394C";
    when 16#1499# => romdata <= X"C8EB7B82";
    when 16#149A# => romdata <= X"8A60C53A";
    when 16#149B# => romdata <= X"2FEC3315";
    when 16#149C# => romdata <= X"BEAEB300";
    when 16#149D# => romdata <= X"45B3E650";
    when 16#149E# => romdata <= X"06C6EBB2";
    when 16#149F# => romdata <= X"3B47A8A0";
    when 16#14A0# => romdata <= X"69EAD45E";
    when 16#14A1# => romdata <= X"32E771B9";
    when 16#14A2# => romdata <= X"C467B435";
    when 16#14A3# => romdata <= X"9EBB681A";
    when 16#14A4# => romdata <= X"B48C891A";
    when 16#14A5# => romdata <= X"BB796544";
    when 16#14A6# => romdata <= X"16917820";
    when 16#14A7# => romdata <= X"3BCC4BC6";
    when 16#14A8# => romdata <= X"B4A278DC";
    when 16#14A9# => romdata <= X"EFACE5E9";
    when 16#14AA# => romdata <= X"385C0593";
    when 16#14AB# => romdata <= X"46A23DCC";
    when 16#14AC# => romdata <= X"A001FC9E";
    when 16#14AD# => romdata <= X"47CFEED4";
    when 16#14AE# => romdata <= X"BCBDD947";
    when 16#14AF# => romdata <= X"B12A3F7E";
    when 16#14B0# => romdata <= X"5FF8B937";
    when 16#14B1# => romdata <= X"2D9497EE";
    when 16#14B2# => romdata <= X"1A508D8B";
    when 16#14B3# => romdata <= X"D3392BF3";
    when 16#14B4# => romdata <= X"CFAD58F0";
    when 16#14B5# => romdata <= X"191B18F6";
    when 16#14B6# => romdata <= X"A300FF9C";
    when 16#14B7# => romdata <= X"B8D914FD";
    when 16#14B8# => romdata <= X"F37B48BF";
    when 16#14B9# => romdata <= X"24C2C5CA";
    when 16#14BA# => romdata <= X"76ABDFCC";
    when 16#14BB# => romdata <= X"F833D51D";
    when 16#14BC# => romdata <= X"48FC90E0";
    when 16#14BD# => romdata <= X"6E7B9729";
    when 16#14BE# => romdata <= X"44BCBAD1";
    when 16#14BF# => romdata <= X"69232A84";
    when 16#14C0# => romdata <= X"29B6100B";
    when 16#14C1# => romdata <= X"A562F7F3";
    when 16#14C2# => romdata <= X"C55A625A";
    when 16#14C3# => romdata <= X"1870A7C7";
    when 16#14C4# => romdata <= X"D7BC9BD4";
    when 16#14C5# => romdata <= X"C4783278";
    when 16#14C6# => romdata <= X"CD95D07F";
    when 16#14C7# => romdata <= X"89E8010E";
    when 16#14C8# => romdata <= X"78876547";
    when 16#14C9# => romdata <= X"F9AEC443";
    when 16#14CA# => romdata <= X"22B0029A";
    when 16#14CB# => romdata <= X"922B2922";
    when 16#14CC# => romdata <= X"634ECCF2";
    when 16#14CD# => romdata <= X"BBB47BF8";
    when 16#14CE# => romdata <= X"7909C494";
    when 16#14CF# => romdata <= X"049550F1";
    when 16#14D0# => romdata <= X"E6D03BB5";
    when 16#14D1# => romdata <= X"354DEA7E";
    when 16#14D2# => romdata <= X"777F499D";
    when 16#14D3# => romdata <= X"2D6239BF";
    when 16#14D4# => romdata <= X"A5C1CFA5";
    when 16#14D5# => romdata <= X"36F8CB16";
    when 16#14D6# => romdata <= X"F4DB9EAD";
    when 16#14D7# => romdata <= X"96F83A4A";
    when 16#14D8# => romdata <= X"D34AE2C6";
    when 16#14D9# => romdata <= X"893ECD69";
    when 16#14DA# => romdata <= X"94C89E7F";
    when 16#14DB# => romdata <= X"4FE426D9";
    when 16#14DC# => romdata <= X"5A18F93B";
    when 16#14DD# => romdata <= X"88CB3579";
    when 16#14DE# => romdata <= X"96B8E5A3";
    when 16#14DF# => romdata <= X"4C43533E";
    when 16#14E0# => romdata <= X"DB1F28A8";
    when 16#14E1# => romdata <= X"162FCBEF";
    when 16#14E2# => romdata <= X"03704FCC";
    when 16#14E3# => romdata <= X"CD80C328";
    when 16#14E4# => romdata <= X"74F345D3";
    when 16#14E5# => romdata <= X"4E81EE81";
    when 16#14E6# => romdata <= X"3DF5CC9B";
    when 16#14E7# => romdata <= X"9C299362";
    when 16#14E8# => romdata <= X"F8443AAB";
    when 16#14E9# => romdata <= X"E91BD0EA";
    when 16#14EA# => romdata <= X"B9746E43";
    when 16#14EB# => romdata <= X"1804B612";
    when 16#14EC# => romdata <= X"9FD32916";
    when 16#14ED# => romdata <= X"303A5703";
    when 16#14EE# => romdata <= X"23FA121F";
    when 16#14EF# => romdata <= X"7AEB2829";
    when 16#14F0# => romdata <= X"F2A50A82";
    when 16#14F1# => romdata <= X"CACCF6D2";
    when 16#14F2# => romdata <= X"73FFBD7A";
    when 16#14F3# => romdata <= X"C6FFC580";
    when 16#14F4# => romdata <= X"7771D216";
    when 16#14F5# => romdata <= X"F50742F7";
    when 16#14F6# => romdata <= X"091946F9";
    when 16#14F7# => romdata <= X"14601159";
    when 16#14F8# => romdata <= X"89C87E8B";
    when 16#14F9# => romdata <= X"BBC8402B";
    when 16#14FA# => romdata <= X"4C8B95C1";
    when 16#14FB# => romdata <= X"02CAB538";
    when 16#14FC# => romdata <= X"43D581FA";
    when 16#14FD# => romdata <= X"9F16C0EC";
    when 16#14FE# => romdata <= X"CE8944E5";
    when 16#14FF# => romdata <= X"FC4BF4C0";
    when 16#1500# => romdata <= X"9D7B1CF0";
    when 16#1501# => romdata <= X"029261D6";
    when 16#1502# => romdata <= X"5AE1F021";
    when 16#1503# => romdata <= X"DAFA81CF";
    when 16#1504# => romdata <= X"1673C9E0";
    when 16#1505# => romdata <= X"B47FF2C3";
    when 16#1506# => romdata <= X"7D1B1AF4";
    when 16#1507# => romdata <= X"6E7A91BC";
    when 16#1508# => romdata <= X"5E529C8F";
    when 16#1509# => romdata <= X"93EE3BC7";
    when 16#150A# => romdata <= X"4E92B274";
    when 16#150B# => romdata <= X"3AAB1EDE";
    when 16#150C# => romdata <= X"16A6523B";
    when 16#150D# => romdata <= X"5B8A591C";
    when 16#150E# => romdata <= X"617C1FD0";
    when 16#150F# => romdata <= X"150E63F3";
    when 16#1510# => romdata <= X"B7EF0494";
    when 16#1511# => romdata <= X"162437B0";
    when 16#1512# => romdata <= X"FD555A83";
    when 16#1513# => romdata <= X"A3BDB519";
    when 16#1514# => romdata <= X"B3BB209E";
    when 16#1515# => romdata <= X"F7924D6B";
    when 16#1516# => romdata <= X"CDE5992B";
    when 16#1517# => romdata <= X"A6248690";
    when 16#1518# => romdata <= X"442E72CD";
    when 16#1519# => romdata <= X"5EB64B4C";
    when 16#151A# => romdata <= X"3D3F7DA3";
    when 16#151B# => romdata <= X"39108A18";
    when 16#151C# => romdata <= X"B61AD88A";
    when 16#151D# => romdata <= X"BE87BB7C";
    when 16#151E# => romdata <= X"85A3A352";
    when 16#151F# => romdata <= X"D7B882FD";
    when 16#1520# => romdata <= X"683B2637";
    when 16#1521# => romdata <= X"A17A2D9C";
    when 16#1522# => romdata <= X"B0B7F414";
    when 16#1523# => romdata <= X"56DCFA66";
    when 16#1524# => romdata <= X"D62913F1";
    when 16#1525# => romdata <= X"45600BAA";
    when 16#1526# => romdata <= X"EEE7EFA5";
    when 16#1527# => romdata <= X"071C3C9E";
    when 16#1528# => romdata <= X"6FDD0A67";
    when 16#1529# => romdata <= X"79A73707";
    when 16#152A# => romdata <= X"1FA69659";
    when 16#152B# => romdata <= X"78CBC897";
    when 16#152C# => romdata <= X"76386B10";
    when 16#152D# => romdata <= X"8DD7216F";
    when 16#152E# => romdata <= X"CE962FA8";
    when 16#152F# => romdata <= X"7A26B29F";
    when 16#1530# => romdata <= X"E0E73230";
    when 16#1531# => romdata <= X"9C0124B0";
    when 16#1532# => romdata <= X"C1E99E56";
    when 16#1533# => romdata <= X"42E5EAE6";
    when 16#1534# => romdata <= X"70005B07";
    when 16#1535# => romdata <= X"8C097D16";
    when 16#1536# => romdata <= X"C58B8923";
    when 16#1537# => romdata <= X"633C18FD";
    when 16#1538# => romdata <= X"B0E8FF8C";
    when 16#1539# => romdata <= X"4610B789";
    when 16#153A# => romdata <= X"387ACB5A";
    when 16#153B# => romdata <= X"2DD0B6AE";
    when 16#153C# => romdata <= X"7E0DF43A";
    when 16#153D# => romdata <= X"6A9E8C3B";
    when 16#153E# => romdata <= X"89C7E5D6";
    when 16#153F# => romdata <= X"28D59759";
    when 16#1540# => romdata <= X"C58D07E0";
    when 16#1541# => romdata <= X"687812AE";
    when 16#1542# => romdata <= X"DAEEDBC6";
    when 16#1543# => romdata <= X"3B4FEE85";
    when 16#1544# => romdata <= X"24D10E4B";
    when 16#1545# => romdata <= X"46769695";
    when 16#1546# => romdata <= X"7E6791C1";
    when 16#1547# => romdata <= X"E94B13CA";
    when 16#1548# => romdata <= X"DCD0ED60";
    when 16#1549# => romdata <= X"752C2DB1";
    when 16#154A# => romdata <= X"B65E035E";
    when 16#154B# => romdata <= X"A72F89FC";
    when 16#154C# => romdata <= X"679138D3";
    when 16#154D# => romdata <= X"609FD2A3";
    when 16#154E# => romdata <= X"0E4DD1A9";
    when 16#154F# => romdata <= X"46418253";
    when 16#1550# => romdata <= X"C67AA69B";
    when 16#1551# => romdata <= X"07EBB95D";
    when 16#1552# => romdata <= X"4973F562";
    when 16#1553# => romdata <= X"CE377343";
    when 16#1554# => romdata <= X"0007A6DB";
    when 16#1555# => romdata <= X"77271D5F";
    when 16#1556# => romdata <= X"2B342CC5";
    when 16#1557# => romdata <= X"E76E1151";
    when 16#1558# => romdata <= X"78F9C7B1";
    when 16#1559# => romdata <= X"600554F5";
    when 16#155A# => romdata <= X"C794961B";
    when 16#155B# => romdata <= X"AE81A5E9";
    when 16#155C# => romdata <= X"B621BA17";
    when 16#155D# => romdata <= X"851008BE";
    when 16#155E# => romdata <= X"D9B556E4";
    when 16#155F# => romdata <= X"61A553FE";
    when 16#1560# => romdata <= X"9BE00A40";
    when 16#1561# => romdata <= X"891750E4";
    when 16#1562# => romdata <= X"EA4B4752";
    when 16#1563# => romdata <= X"16283B53";
    when 16#1564# => romdata <= X"0CB8D479";
    when 16#1565# => romdata <= X"DC70B026";
    when 16#1566# => romdata <= X"E0788922";
    when 16#1567# => romdata <= X"9F601755";
    when 16#1568# => romdata <= X"2AB9E01E";
    when 16#1569# => romdata <= X"DE6703FD";
    when 16#156A# => romdata <= X"1E2D59AF";
    when 16#156B# => romdata <= X"0B71E0F1";
    when 16#156C# => romdata <= X"DC9A42AC";
    when 16#156D# => romdata <= X"C5823324";
    when 16#156E# => romdata <= X"BEFC52CA";
    when 16#156F# => romdata <= X"0DCD25FE";
    when 16#1570# => romdata <= X"8B10C999";
    when 16#1571# => romdata <= X"152AA367";
    when 16#1572# => romdata <= X"6A30602D";
    when 16#1573# => romdata <= X"3506F787";
    when 16#1574# => romdata <= X"51477033";
    when 16#1575# => romdata <= X"DB7AB1A2";
    when 16#1576# => romdata <= X"EDC21A6F";
    when 16#1577# => romdata <= X"E51273B6";
    when 16#1578# => romdata <= X"B2890088";
    when 16#1579# => romdata <= X"703CEFE7";
    when 16#157A# => romdata <= X"4F9EA898";
    when 16#157B# => romdata <= X"81896E5B";
    when 16#157C# => romdata <= X"E124B1FC";
    when 16#157D# => romdata <= X"9430B92F";
    when 16#157E# => romdata <= X"0C0568F5";
    when 16#157F# => romdata <= X"A068A800";
    when 16#1580# => romdata <= X"F23088E3";
    when 16#1581# => romdata <= X"EAA0A6BA";
    when 16#1582# => romdata <= X"04D0633A";
    when 16#1583# => romdata <= X"AFE85203";
    when 16#1584# => romdata <= X"E8B18292";
    when 16#1585# => romdata <= X"23FA6B73";
    when 16#1586# => romdata <= X"0F6DEE67";
    when 16#1587# => romdata <= X"99B521F2";
    when 16#1588# => romdata <= X"E8323B87";
    when 16#1589# => romdata <= X"93D0F7F2";
    when 16#158A# => romdata <= X"BB9305B3";
    when 16#158B# => romdata <= X"EF4F5B4F";
    when 16#158C# => romdata <= X"1CB82283";
    when 16#158D# => romdata <= X"6E4D92C8";
    when 16#158E# => romdata <= X"E4928A85";
    when 16#158F# => romdata <= X"1BCE6883";
    when 16#1590# => romdata <= X"29DECA6F";
    when 16#1591# => romdata <= X"7285DCC8";
    when 16#1592# => romdata <= X"5195E5BD";
    when 16#1593# => romdata <= X"A3B503B8";
    when 16#1594# => romdata <= X"AEE6F1CD";
    when 16#1595# => romdata <= X"7FBB1584";
    when 16#1596# => romdata <= X"44E7DE8B";
    when 16#1597# => romdata <= X"F6A9A3CD";
    when 16#1598# => romdata <= X"A3117877";
    when 16#1599# => romdata <= X"55A827BC";
    when 16#159A# => romdata <= X"AD3DA562";
    when 16#159B# => romdata <= X"1908EA91";
    when 16#159C# => romdata <= X"3C0316B9";
    when 16#159D# => romdata <= X"B52BFB07";
    when 16#159E# => romdata <= X"ADADEFF1";
    when 16#159F# => romdata <= X"7D3766BB";
    when 16#15A0# => romdata <= X"450DD713";
    when 16#15A1# => romdata <= X"28A0353B";
    when 16#15A2# => romdata <= X"09DC24DE";
    when 16#15A3# => romdata <= X"93CF83A2";
    when 16#15A4# => romdata <= X"E5F98BA9";
    when 16#15A5# => romdata <= X"D612187B";
    when 16#15A6# => romdata <= X"601157D6";
    when 16#15A7# => romdata <= X"B140E675";
    when 16#15A8# => romdata <= X"228B58C9";
    when 16#15A9# => romdata <= X"398618C3";
    when 16#15AA# => romdata <= X"BF0D11A2";
    when 16#15AB# => romdata <= X"26E48936";
    when 16#15AC# => romdata <= X"6102B9C3";
    when 16#15AD# => romdata <= X"5A916653";
    when 16#15AE# => romdata <= X"F0DB3671";
    when 16#15AF# => romdata <= X"1ACBA5F3";
    when 16#15B0# => romdata <= X"2B327F57";
    when 16#15B1# => romdata <= X"89F3EF48";
    when 16#15B2# => romdata <= X"A338E467";
    when 16#15B3# => romdata <= X"6F4BC2C6";
    when 16#15B4# => romdata <= X"A1308597";
    when 16#15B5# => romdata <= X"171903D2";
    when 16#15B6# => romdata <= X"AA299CE7";
    when 16#15B7# => romdata <= X"E523C2AB";
    when 16#15B8# => romdata <= X"E4B15AA4";
    when 16#15B9# => romdata <= X"FC489541";
    when 16#15BA# => romdata <= X"87E00975";
    when 16#15BB# => romdata <= X"83EB0994";
    when 16#15BC# => romdata <= X"19047244";
    when 16#15BD# => romdata <= X"B4931326";
    when 16#15BE# => romdata <= X"E5923B63";
    when 16#15BF# => romdata <= X"13DE0842";
    when 16#15C0# => romdata <= X"3DB00866";
    when 16#15C1# => romdata <= X"374ABBF5";
    when 16#15C2# => romdata <= X"C31A0054";
    when 16#15C3# => romdata <= X"2CB97CDF";
    when 16#15C4# => romdata <= X"B8F71046";
    when 16#15C5# => romdata <= X"AA2A6DBF";
    when 16#15C6# => romdata <= X"D7E1A71C";
    when 16#15C7# => romdata <= X"068ED70E";
    when 16#15C8# => romdata <= X"8D7C3268";
    when 16#15C9# => romdata <= X"EA3E0EEF";
    when 16#15CA# => romdata <= X"2262BD79";
    when 16#15CB# => romdata <= X"91B6C59F";
    when 16#15CC# => romdata <= X"F471F73A";
    when 16#15CD# => romdata <= X"4E85F4FA";
    when 16#15CE# => romdata <= X"015E164F";
    when 16#15CF# => romdata <= X"9C15FE0A";
    when 16#15D0# => romdata <= X"A5F4772B";
    when 16#15D1# => romdata <= X"F2D62B26";
    when 16#15D2# => romdata <= X"D3EAA25C";
    when 16#15D3# => romdata <= X"E83EAEC5";
    when 16#15D4# => romdata <= X"EB3577CA";
    when 16#15D5# => romdata <= X"83A68168";
    when 16#15D6# => romdata <= X"FB64C40A";
    when 16#15D7# => romdata <= X"7A155905";
    when 16#15D8# => romdata <= X"CBA6E641";
    when 16#15D9# => romdata <= X"59E55EBC";
    when 16#15DA# => romdata <= X"928D125E";
    when 16#15DB# => romdata <= X"55165C63";
    when 16#15DC# => romdata <= X"9F545B00";
    when 16#15DD# => romdata <= X"71EE3CF1";
    when 16#15DE# => romdata <= X"A3F58B49";
    when 16#15DF# => romdata <= X"94BB4BF5";
    when 16#15E0# => romdata <= X"0C2B24F2";
    when 16#15E1# => romdata <= X"E06E4ADC";
    when 16#15E2# => romdata <= X"90BC1C09";
    when 16#15E3# => romdata <= X"54A257D8";
    when 16#15E4# => romdata <= X"8444347A";
    when 16#15E5# => romdata <= X"AECF136C";
    when 16#15E6# => romdata <= X"15242633";
    when 16#15E7# => romdata <= X"463DCF98";
    when 16#15E8# => romdata <= X"4BB67366";
    when 16#15E9# => romdata <= X"66E38F1A";
    when 16#15EA# => romdata <= X"45150B1B";
    when 16#15EB# => romdata <= X"7D1C31DE";
    when 16#15EC# => romdata <= X"06EB9C2F";
    when 16#15ED# => romdata <= X"4097E9D9";
    when 16#15EE# => romdata <= X"B4D21EBC";
    when 16#15EF# => romdata <= X"9F3A9180";
    when 16#15F0# => romdata <= X"00DE2449";
    when 16#15F1# => romdata <= X"DCB3F5FD";
    when 16#15F2# => romdata <= X"DC3C773A";
    when 16#15F3# => romdata <= X"645DF560";
    when 16#15F4# => romdata <= X"F7E013E8";
    when 16#15F5# => romdata <= X"47E2356D";
    when 16#15F6# => romdata <= X"33EFF1E2";
    when 16#15F7# => romdata <= X"15782638";
    when 16#15F8# => romdata <= X"F58034B0";
    when 16#15F9# => romdata <= X"9F4739F9";
    when 16#15FA# => romdata <= X"8915BFB0";
    when 16#15FB# => romdata <= X"B1DC1246";
    when 16#15FC# => romdata <= X"81492F58";
    when 16#15FD# => romdata <= X"021670D0";
    when 16#15FE# => romdata <= X"3CBF5E8F";
    when 16#15FF# => romdata <= X"962351E0";
    when 16#1600# => romdata <= X"EB07F9ED";
    when 16#1601# => romdata <= X"F03596AD";
    when 16#1602# => romdata <= X"C2A3B7EB";
    when 16#1603# => romdata <= X"6DB1CFC9";
    when 16#1604# => romdata <= X"11E9A4C4";
    when 16#1605# => romdata <= X"2336A573";
    when 16#1606# => romdata <= X"09F7B6C3";
    when 16#1607# => romdata <= X"389282E5";
    when 16#1608# => romdata <= X"57D94BCC";
    when 16#1609# => romdata <= X"71827D7C";
    when 16#160A# => romdata <= X"5737B1C5";
    when 16#160B# => romdata <= X"30D2A087";
    when 16#160C# => romdata <= X"E3F50724";
    when 16#160D# => romdata <= X"2F3DA5BD";
    when 16#160E# => romdata <= X"1BBCA4DF";
    when 16#160F# => romdata <= X"8B78BEEC";
    when 16#1610# => romdata <= X"1DBF7EBB";
    when 16#1611# => romdata <= X"2EA1CF1D";
    when 16#1612# => romdata <= X"FA79E607";
    when 16#1613# => romdata <= X"85BAFA23";
    when 16#1614# => romdata <= X"658490C9";
    when 16#1615# => romdata <= X"A64AC61C";
    when 16#1616# => romdata <= X"45779DFA";
    when 16#1617# => romdata <= X"FC6C55CB";
    when 16#1618# => romdata <= X"5C9FE457";
    when 16#1619# => romdata <= X"BF47E45A";
    when 16#161A# => romdata <= X"3FEF092E";
    when 16#161B# => romdata <= X"178ED449";
    when 16#161C# => romdata <= X"5C0357B4";
    when 16#161D# => romdata <= X"59E95AAC";
    when 16#161E# => romdata <= X"82132FF1";
    when 16#161F# => romdata <= X"C8044F4E";
    when 16#1620# => romdata <= X"C84EB882";
    when 16#1621# => romdata <= X"DC195D9C";
    when 16#1622# => romdata <= X"E996B1CC";
    when 16#1623# => romdata <= X"F523098E";
    when 16#1624# => romdata <= X"9E1A57C3";
    when 16#1625# => romdata <= X"7C2E2D0A";
    when 16#1626# => romdata <= X"CB0EAA34";
    when 16#1627# => romdata <= X"B0B56FE5";
    when 16#1628# => romdata <= X"A0747130";
    when 16#1629# => romdata <= X"B1E75AA9";
    when 16#162A# => romdata <= X"23F6F94C";
    when 16#162B# => romdata <= X"0D024A7F";
    when 16#162C# => romdata <= X"CD22E7A4";
    when 16#162D# => romdata <= X"ED8B2019";
    when 16#162E# => romdata <= X"66C417AE";
    when 16#162F# => romdata <= X"86442076";
    when 16#1630# => romdata <= X"7AB3223B";
    when 16#1631# => romdata <= X"FF56C64D";
    when 16#1632# => romdata <= X"4F8F557D";
    when 16#1633# => romdata <= X"D950F7C5";
    when 16#1634# => romdata <= X"0D9A39AB";
    when 16#1635# => romdata <= X"2C742CE6";
    when 16#1636# => romdata <= X"86C8F92B";
    when 16#1637# => romdata <= X"35711904";
    when 16#1638# => romdata <= X"C600A9D4";
    when 16#1639# => romdata <= X"D3DD83F3";
    when 16#163A# => romdata <= X"DF1ED7DB";
    when 16#163B# => romdata <= X"8042C76B";
    when 16#163C# => romdata <= X"0B7D5D9B";
    when 16#163D# => romdata <= X"CD6E0B55";
    when 16#163E# => romdata <= X"24184BF9";
    when 16#163F# => romdata <= X"9D8D0B4F";
    when 16#1640# => romdata <= X"14967FA4";
    when 16#1641# => romdata <= X"8A93A2F4";
    when 16#1642# => romdata <= X"4E2275ED";
    when 16#1643# => romdata <= X"7E59F399";
    when 16#1644# => romdata <= X"1EFB0CBF";
    when 16#1645# => romdata <= X"2E26AC1F";
    when 16#1646# => romdata <= X"8D9A41AA";
    when 16#1647# => romdata <= X"E4563179";
    when 16#1648# => romdata <= X"254BA370";
    when 16#1649# => romdata <= X"28867E68";
    when 16#164A# => romdata <= X"C8179454";
    when 16#164B# => romdata <= X"B8B71FAB";
    when 16#164C# => romdata <= X"49DBD1F8";
    when 16#164D# => romdata <= X"89104CFB";
    when 16#164E# => romdata <= X"64C81211";
    when 16#164F# => romdata <= X"51364BDB";
    when 16#1650# => romdata <= X"64BAF854";
    when 16#1651# => romdata <= X"B0DA22B8";
    when 16#1652# => romdata <= X"620BD7EE";
    when 16#1653# => romdata <= X"3D4302A8";
    when 16#1654# => romdata <= X"8A115F8B";
    when 16#1655# => romdata <= X"FBA649CA";
    when 16#1656# => romdata <= X"A9EE7EF5";
    when 16#1657# => romdata <= X"BC95CFAB";
    when 16#1658# => romdata <= X"26503A9D";
    when 16#1659# => romdata <= X"26033370";
    when 16#165A# => romdata <= X"A4EF3CB8";
    when 16#165B# => romdata <= X"A5D094C6";
    when 16#165C# => romdata <= X"3305A833";
    when 16#165D# => romdata <= X"387B4F83";
    when 16#165E# => romdata <= X"71C6FE19";
    when 16#165F# => romdata <= X"87514BB4";
    when 16#1660# => romdata <= X"58C571E6";
    when 16#1661# => romdata <= X"CB5DF5FC";
    when 16#1662# => romdata <= X"90063165";
    when 16#1663# => romdata <= X"2D3FA444";
    when 16#1664# => romdata <= X"4F8F1F03";
    when 16#1665# => romdata <= X"12204340";
    when 16#1666# => romdata <= X"FDB2092F";
    when 16#1667# => romdata <= X"709FDC51";
    when 16#1668# => romdata <= X"D2680753";
    when 16#1669# => romdata <= X"131ABC33";
    when 16#166A# => romdata <= X"712B4F10";
    when 16#166B# => romdata <= X"67EA1CC8";
    when 16#166C# => romdata <= X"7C40B281";
    when 16#166D# => romdata <= X"E69209ED";
    when 16#166E# => romdata <= X"EC42C22A";
    when 16#166F# => romdata <= X"88950E9C";
    when 16#1670# => romdata <= X"1CE8130D";
    when 16#1671# => romdata <= X"A9291897";
    when 16#1672# => romdata <= X"BF2D8D1D";
    when 16#1673# => romdata <= X"10691174";
    when 16#1674# => romdata <= X"3E7A9DA3";
    when 16#1675# => romdata <= X"6220FA90";
    when 16#1676# => romdata <= X"A02A34EB";
    when 16#1677# => romdata <= X"0B285432";
    when 16#1678# => romdata <= X"17839374";
    when 16#1679# => romdata <= X"EBE79F40";
    when 16#167A# => romdata <= X"B3B61223";
    when 16#167B# => romdata <= X"6C902E4C";
    when 16#167C# => romdata <= X"D05CE2E1";
    when 16#167D# => romdata <= X"C07F3DA1";
    when 16#167E# => romdata <= X"0E2AEE8E";
    when 16#167F# => romdata <= X"387494E0";
    when 16#1680# => romdata <= X"E9D537A8";
    when 16#1681# => romdata <= X"21DEDE52";
    when 16#1682# => romdata <= X"6B441BA4";
    when 16#1683# => romdata <= X"25278577";
    when 16#1684# => romdata <= X"9B54DE76";
    when 16#1685# => romdata <= X"F82747F8";
    when 16#1686# => romdata <= X"607B8952";
    when 16#1687# => romdata <= X"DF990F26";
    when 16#1688# => romdata <= X"8C039CC7";
    when 16#1689# => romdata <= X"92883B1C";
    when 16#168A# => romdata <= X"76C297D8";
    when 16#168B# => romdata <= X"1C6C0CF1";
    when 16#168C# => romdata <= X"7DA8BA2C";
    when 16#168D# => romdata <= X"71110B16";
    when 16#168E# => romdata <= X"74172872";
    when 16#168F# => romdata <= X"5839D33B";
    when 16#1690# => romdata <= X"5942BC0A";
    when 16#1691# => romdata <= X"5614A365";
    when 16#1692# => romdata <= X"0675FDA5";
    when 16#1693# => romdata <= X"D70F2915";
    when 16#1694# => romdata <= X"4A429A42";
    when 16#1695# => romdata <= X"819D6EDE";
    when 16#1696# => romdata <= X"324C6459";
    when 16#1697# => romdata <= X"6F93E84C";
    when 16#1698# => romdata <= X"C9B2C9DA";
    when 16#1699# => romdata <= X"3717AA6D";
    when 16#169A# => romdata <= X"FFCD03B7";
    when 16#169B# => romdata <= X"5AC96543";
    when 16#169C# => romdata <= X"020A9F20";
    when 16#169D# => romdata <= X"24620353";
    when 16#169E# => romdata <= X"E1364E43";
    when 16#169F# => romdata <= X"20FD4493";
    when 16#16A0# => romdata <= X"3799FFF0";
    when 16#16A1# => romdata <= X"83E73F5D";
    when 16#16A2# => romdata <= X"20B83BF7";
    when 16#16A3# => romdata <= X"7EC22479";
    when 16#16A4# => romdata <= X"64ECE442";
    when 16#16A5# => romdata <= X"C3213DE9";
    when 16#16A6# => romdata <= X"9026F8FA";
    when 16#16A7# => romdata <= X"F0E96302";
    when 16#16A8# => romdata <= X"EC60067E";
    when 16#16A9# => romdata <= X"A38C5CA0";
    when 16#16AA# => romdata <= X"CD989475";
    when 16#16AB# => romdata <= X"205FA388";
    when 16#16AC# => romdata <= X"69E349FC";
    when 16#16AD# => romdata <= X"7F79EB81";
    when 16#16AE# => romdata <= X"F8457CA3";
    when 16#16AF# => romdata <= X"D1A875A8";
    when 16#16B0# => romdata <= X"D166C96E";
    when 16#16B1# => romdata <= X"BAF1F39C";
    when 16#16B2# => romdata <= X"88815E22";
    when 16#16B3# => romdata <= X"58EA1A14";
    when 16#16B4# => romdata <= X"943298DA";
    when 16#16B5# => romdata <= X"39EB9B73";
    when 16#16B6# => romdata <= X"8AAA4E00";
    when 16#16B7# => romdata <= X"35F9567A";
    when 16#16B8# => romdata <= X"0A9D5727";
    when 16#16B9# => romdata <= X"85594496";
    when 16#16BA# => romdata <= X"316D56EB";
    when 16#16BB# => romdata <= X"3D39E1F3";
    when 16#16BC# => romdata <= X"F243D4F1";
    when 16#16BD# => romdata <= X"6111E194";
    when 16#16BE# => romdata <= X"FC537A63";
    when 16#16BF# => romdata <= X"5FAEB2FB";
    when 16#16C0# => romdata <= X"4401CAA9";
    when 16#16C1# => romdata <= X"EE0091CF";
    when 16#16C2# => romdata <= X"3CB28B36";
    when 16#16C3# => romdata <= X"6CB5446A";
    when 16#16C4# => romdata <= X"6D3B10AB";
    when 16#16C5# => romdata <= X"86B4B1A0";
    when 16#16C6# => romdata <= X"714D107F";
    when 16#16C7# => romdata <= X"CCBBD50E";
    when 16#16C8# => romdata <= X"AE520D56";
    when 16#16C9# => romdata <= X"A1161E03";
    when 16#16CA# => romdata <= X"849192F5";
    when 16#16CB# => romdata <= X"096346FB";
    when 16#16CC# => romdata <= X"E5150B6D";
    when 16#16CD# => romdata <= X"04025A56";
    when 16#16CE# => romdata <= X"4A43A3D2";
    when 16#16CF# => romdata <= X"2BD4B7E1";
    when 16#16D0# => romdata <= X"0DD4061C";
    when 16#16D1# => romdata <= X"E20FA2EC";
    when 16#16D2# => romdata <= X"DD36F66B";
    when 16#16D3# => romdata <= X"AAD7EA96";
    when 16#16D4# => romdata <= X"CDBAA0F0";
    when 16#16D5# => romdata <= X"63B81470";
    when 16#16D6# => romdata <= X"7718F472";
    when 16#16D7# => romdata <= X"78F8570F";
    when 16#16D8# => romdata <= X"77F3B157";
    when 16#16D9# => romdata <= X"99D0E354";
    when 16#16DA# => romdata <= X"CCA50DAA";
    when 16#16DB# => romdata <= X"38C31C74";
    when 16#16DC# => romdata <= X"6B174822";
    when 16#16DD# => romdata <= X"97D9C089";
    when 16#16DE# => romdata <= X"FF379454";
    when 16#16DF# => romdata <= X"FCCCB873";
    when 16#16E0# => romdata <= X"0D89B146";
    when 16#16E1# => romdata <= X"2AD95426";
    when 16#16E2# => romdata <= X"370AC37D";
    when 16#16E3# => romdata <= X"E50B775B";
    when 16#16E4# => romdata <= X"952663B9";
    when 16#16E5# => romdata <= X"7AFBC403";
    when 16#16E6# => romdata <= X"F6F729BB";
    when 16#16E7# => romdata <= X"9CC1D21D";
    when 16#16E8# => romdata <= X"D89EE78A";
    when 16#16E9# => romdata <= X"F09DF855";
    when 16#16EA# => romdata <= X"8F7E68B3";
    when 16#16EB# => romdata <= X"711A7D90";
    when 16#16EC# => romdata <= X"75DD4754";
    when 16#16ED# => romdata <= X"174802F5";
    when 16#16EE# => romdata <= X"2CB9683F";
    when 16#16EF# => romdata <= X"FE746471";
    when 16#16F0# => romdata <= X"C7E543FF";
    when 16#16F1# => romdata <= X"388D0243";
    when 16#16F2# => romdata <= X"27D1866C";
    when 16#16F3# => romdata <= X"C5CA6775";
    when 16#16F4# => romdata <= X"C58A14D7";
    when 16#16F5# => romdata <= X"0A3ECCD3";
    when 16#16F6# => romdata <= X"EFAB52F9";
    when 16#16F7# => romdata <= X"AE6CCE14";
    when 16#16F8# => romdata <= X"6766A841";
    when 16#16F9# => romdata <= X"9FB546E3";
    when 16#16FA# => romdata <= X"9EB604F4";
    when 16#16FB# => romdata <= X"3B15AB88";
    when 16#16FC# => romdata <= X"C72741F8";
    when 16#16FD# => romdata <= X"C7D0A7FE";
    when 16#16FE# => romdata <= X"2F462D36";
    when 16#16FF# => romdata <= X"0676D6E0";
    when 16#1700# => romdata <= X"D79D9162";
    when 16#1701# => romdata <= X"41BBE52B";
    when 16#1702# => romdata <= X"61BE8210";
    when 16#1703# => romdata <= X"A02543F7";
    when 16#1704# => romdata <= X"5A47032E";
    when 16#1705# => romdata <= X"9C0CC128";
    when 16#1706# => romdata <= X"524A675E";
    when 16#1707# => romdata <= X"94D8F79A";
    when 16#1708# => romdata <= X"69B6842B";
    when 16#1709# => romdata <= X"0C5CFF5C";
    when 16#170A# => romdata <= X"1AC98D20";
    when 16#170B# => romdata <= X"85299BDB";
    when 16#170C# => romdata <= X"AEA67A41";
    when 16#170D# => romdata <= X"C724CA36";
    when 16#170E# => romdata <= X"B6275A80";
    when 16#170F# => romdata <= X"D377DC3A";
    when 16#1710# => romdata <= X"6EB4C8D0";
    when 16#1711# => romdata <= X"B6B88241";
    when 16#1712# => romdata <= X"334A9530";
    when 16#1713# => romdata <= X"0B53FFB5";
    when 16#1714# => romdata <= X"46163D28";
    when 16#1715# => romdata <= X"89D7C85F";
    when 16#1716# => romdata <= X"1D139792";
    when 16#1717# => romdata <= X"4F126DA7";
    when 16#1718# => romdata <= X"6085BEF1";
    when 16#1719# => romdata <= X"31A65C7D";
    when 16#171A# => romdata <= X"DF60DDF4";
    when 16#171B# => romdata <= X"086BD33B";
    when 16#171C# => romdata <= X"44D25025";
    when 16#171D# => romdata <= X"D689FF41";
    when 16#171E# => romdata <= X"E0C256EA";
    when 16#171F# => romdata <= X"12F4353D";
    when 16#1720# => romdata <= X"9E722EE3";
    when 16#1721# => romdata <= X"7907AA8B";
    when 16#1722# => romdata <= X"ED0A5A60";
    when 16#1723# => romdata <= X"6333A031";
    when 16#1724# => romdata <= X"AC6B9A16";
    when 16#1725# => romdata <= X"61425091";
    when 16#1726# => romdata <= X"6759B72F";
    when 16#1727# => romdata <= X"E6C1828B";
    when 16#1728# => romdata <= X"C6C1966C";
    when 16#1729# => romdata <= X"9EBCD514";
    when 16#172A# => romdata <= X"13A77F41";
    when 16#172B# => romdata <= X"F808BCA2";
    when 16#172C# => romdata <= X"534AC49D";
    when 16#172D# => romdata <= X"B1D32D37";
    when 16#172E# => romdata <= X"878DF5CC";
    when 16#172F# => romdata <= X"0BEFCC09";
    when 16#1730# => romdata <= X"9C56CAF5";
    when 16#1731# => romdata <= X"0D8B92E7";
    when 16#1732# => romdata <= X"CE616AA0";
    when 16#1733# => romdata <= X"26EA1D81";
    when 16#1734# => romdata <= X"DC7ABC17";
    when 16#1735# => romdata <= X"C4705F9B";
    when 16#1736# => romdata <= X"57A0F99F";
    when 16#1737# => romdata <= X"A749F30F";
    when 16#1738# => romdata <= X"93DFA982";
    when 16#1739# => romdata <= X"A083EAE6";
    when 16#173A# => romdata <= X"582C8461";
    when 16#173B# => romdata <= X"A11ABA74";
    when 16#173C# => romdata <= X"B11663ED";
    when 16#173D# => romdata <= X"7D66EB4F";
    when 16#173E# => romdata <= X"8DE14F09";
    when 16#173F# => romdata <= X"0EB1CA6D";
    when 16#1740# => romdata <= X"8D81CB6B";
    when 16#1741# => romdata <= X"063A391F";
    when 16#1742# => romdata <= X"D354DCEA";
    when 16#1743# => romdata <= X"F7DB71C2";
    when 16#1744# => romdata <= X"77D0E92B";
    when 16#1745# => romdata <= X"4B463873";
    when 16#1746# => romdata <= X"DCBEFFB6";
    when 16#1747# => romdata <= X"98BDCA17";
    when 16#1748# => romdata <= X"F80845EF";
    when 16#1749# => romdata <= X"D5F0FF15";
    when 16#174A# => romdata <= X"0ADDC9D7";
    when 16#174B# => romdata <= X"797E21E4";
    when 16#174C# => romdata <= X"279B54BD";
    when 16#174D# => romdata <= X"D4B7C9D4";
    when 16#174E# => romdata <= X"03D9FA61";
    when 16#174F# => romdata <= X"01604B79";
    when 16#1750# => romdata <= X"AC377780";
    when 16#1751# => romdata <= X"A5461499";
    when 16#1752# => romdata <= X"71408294";
    when 16#1753# => romdata <= X"2313CF74";
    when 16#1754# => romdata <= X"AD1147CD";
    when 16#1755# => romdata <= X"10571A31";
    when 16#1756# => romdata <= X"D82871B6";
    when 16#1757# => romdata <= X"B3A055D5";
    when 16#1758# => romdata <= X"0C6CDA4B";
    when 16#1759# => romdata <= X"DDF3871F";
    when 16#175A# => romdata <= X"41EFDAEB";
    when 16#175B# => romdata <= X"E8ABB995";
    when 16#175C# => romdata <= X"344DB636";
    when 16#175D# => romdata <= X"6E35C6E5";
    when 16#175E# => romdata <= X"06907AD7";
    when 16#175F# => romdata <= X"FC76632F";
    when 16#1760# => romdata <= X"99124A58";
    when 16#1761# => romdata <= X"A32C8636";
    when 16#1762# => romdata <= X"0FD6DDBF";
    when 16#1763# => romdata <= X"50324D86";
    when 16#1764# => romdata <= X"694518AC";
    when 16#1765# => romdata <= X"44F1FA19";
    when 16#1766# => romdata <= X"662C0EF0";
    when 16#1767# => romdata <= X"C0860811";
    when 16#1768# => romdata <= X"B5B976A9";
    when 16#1769# => romdata <= X"6EC2A144";
    when 16#176A# => romdata <= X"9E53A7E4";
    when 16#176B# => romdata <= X"A07923E9";
    when 16#176C# => romdata <= X"F85794F2";
    when 16#176D# => romdata <= X"28E441D9";
    when 16#176E# => romdata <= X"2903922E";
    when 16#176F# => romdata <= X"5783F2FA";
    when 16#1770# => romdata <= X"21C67725";
    when 16#1771# => romdata <= X"1B6B8DB0";
    when 16#1772# => romdata <= X"2AC2E242";
    when 16#1773# => romdata <= X"C0C8652E";
    when 16#1774# => romdata <= X"0C17C9E3";
    when 16#1775# => romdata <= X"858E52DE";
    when 16#1776# => romdata <= X"78DC712B";
    when 16#1777# => romdata <= X"2DD5D2AF";
    when 16#1778# => romdata <= X"9A42DB2E";
    when 16#1779# => romdata <= X"2BEB3FB6";
    when 16#177A# => romdata <= X"E0FFF13D";
    when 16#177B# => romdata <= X"B9A1E02C";
    when 16#177C# => romdata <= X"8F84FCEF";
    when 16#177D# => romdata <= X"3F7C4D2D";
    when 16#177E# => romdata <= X"DC09F2A2";
    when 16#177F# => romdata <= X"813E8C20";
    when 16#1780# => romdata <= X"F8E2DACD";
    when 16#1781# => romdata <= X"D88277D4";
    when 16#1782# => romdata <= X"82951555";
    when 16#1783# => romdata <= X"C657B3E3";
    when 16#1784# => romdata <= X"C5DB79E5";
    when 16#1785# => romdata <= X"A43500F7";
    when 16#1786# => romdata <= X"A2C8B30C";
    when 16#1787# => romdata <= X"854DBE61";
    when 16#1788# => romdata <= X"1FAC1087";
    when 16#1789# => romdata <= X"FA03D439";
    when 16#178A# => romdata <= X"AC4635D3";
    when 16#178B# => romdata <= X"9211E234";
    when 16#178C# => romdata <= X"B82A9124";
    when 16#178D# => romdata <= X"8DEE5D4F";
    when 16#178E# => romdata <= X"E67A02D5";
    when 16#178F# => romdata <= X"AE25C676";
    when 16#1790# => romdata <= X"E64C4843";
    when 16#1791# => romdata <= X"E419EBB3";
    when 16#1792# => romdata <= X"C4D81FB6";
    when 16#1793# => romdata <= X"06B9CA08";
    when 16#1794# => romdata <= X"36F8207C";
    when 16#1795# => romdata <= X"D19D106C";
    when 16#1796# => romdata <= X"0E287EFD";
    when 16#1797# => romdata <= X"8F8DB5C1";
    when 16#1798# => romdata <= X"A3A22886";
    when 16#1799# => romdata <= X"C2765FED";
    when 16#179A# => romdata <= X"26B51891";
    when 16#179B# => romdata <= X"53657B7C";
    when 16#179C# => romdata <= X"47D5590F";
    when 16#179D# => romdata <= X"11C63400";
    when 16#179E# => romdata <= X"67B80066";
    when 16#179F# => romdata <= X"9B05A084";
    when 16#17A0# => romdata <= X"9BCD2005";
    when 16#17A1# => romdata <= X"DFEE6DF9";
    when 16#17A2# => romdata <= X"5833C9E9";
    when 16#17A3# => romdata <= X"4328D72F";
    when 16#17A4# => romdata <= X"931D69CF";
    when 16#17A5# => romdata <= X"BB2BDA81";
    when 16#17A6# => romdata <= X"AC83DD66";
    when 16#17A7# => romdata <= X"0B3B17D2";
    when 16#17A8# => romdata <= X"BA402349";
    when 16#17A9# => romdata <= X"1DED324F";
    when 16#17AA# => romdata <= X"C4F22510";
    when 16#17AB# => romdata <= X"ECA4A519";
    when 16#17AC# => romdata <= X"4B1245F4";
    when 16#17AD# => romdata <= X"F3FE334D";
    when 16#17AE# => romdata <= X"A9C1E6BF";
    when 16#17AF# => romdata <= X"83A3FB30";
    when 16#17B0# => romdata <= X"897BE54C";
    when 16#17B1# => romdata <= X"688D2A7C";
    when 16#17B2# => romdata <= X"5845F425";
    when 16#17B3# => romdata <= X"866F25DD";
    when 16#17B4# => romdata <= X"0A9852BA";
    when 16#17B5# => romdata <= X"6DAAF843";
    when 16#17B6# => romdata <= X"7DD80BCC";
    when 16#17B7# => romdata <= X"72B3E258";
    when 16#17B8# => romdata <= X"A906DE07";
    when 16#17B9# => romdata <= X"9A2D33EC";
    when 16#17BA# => romdata <= X"5C5F6927";
    when 16#17BB# => romdata <= X"503BA131";
    when 16#17BC# => romdata <= X"58305DFF";
    when 16#17BD# => romdata <= X"D3F86345";
    when 16#17BE# => romdata <= X"52439415";
    when 16#17BF# => romdata <= X"1AA557D6";
    when 16#17C0# => romdata <= X"242060F2";
    when 16#17C1# => romdata <= X"76BB6BB2";
    when 16#17C2# => romdata <= X"5586F632";
    when 16#17C3# => romdata <= X"942ACF5E";
    when 16#17C4# => romdata <= X"0883CD3F";
    when 16#17C5# => romdata <= X"8393688F";
    when 16#17C6# => romdata <= X"360323A0";
    when 16#17C7# => romdata <= X"00B82BD8";
    when 16#17C8# => romdata <= X"9414E9C8";
    when 16#17C9# => romdata <= X"07994B02";
    when 16#17CA# => romdata <= X"34D730BC";
    when 16#17CB# => romdata <= X"6D7CD0A2";
    when 16#17CC# => romdata <= X"BF75D9F5";
    when 16#17CD# => romdata <= X"10786E83";
    when 16#17CE# => romdata <= X"EE98D4CA";
    when 16#17CF# => romdata <= X"CF20EFF8";
    when 16#17D0# => romdata <= X"6EE9C38B";
    when 16#17D1# => romdata <= X"8D52455D";
    when 16#17D2# => romdata <= X"8A694B68";
    when 16#17D3# => romdata <= X"9F0D9A63";
    when 16#17D4# => romdata <= X"2E7A6AC6";
    when 16#17D5# => romdata <= X"675E190A";
    when 16#17D6# => romdata <= X"12ADD716";
    when 16#17D7# => romdata <= X"D2C63226";
    when 16#17D8# => romdata <= X"57B878FA";
    when 16#17D9# => romdata <= X"97267C1B";
    when 16#17DA# => romdata <= X"A4631584";
    when 16#17DB# => romdata <= X"356768EB";
    when 16#17DC# => romdata <= X"BD1F13FD";
    when 16#17DD# => romdata <= X"2F37EBDC";
    when 16#17DE# => romdata <= X"D1DF96FB";
    when 16#17DF# => romdata <= X"943942E8";
    when 16#17E0# => romdata <= X"A5188666";
    when 16#17E1# => romdata <= X"235B455B";
    when 16#17E2# => romdata <= X"E2F770C9";
    when 16#17E3# => romdata <= X"759A8F07";
    when 16#17E4# => romdata <= X"0971CBA4";
    when 16#17E5# => romdata <= X"9789744F";
    when 16#17E6# => romdata <= X"D2F64DC4";
    when 16#17E7# => romdata <= X"DC6E003B";
    when 16#17E8# => romdata <= X"3F9BEC76";
    when 16#17E9# => romdata <= X"17C7EEDF";
    when 16#17EA# => romdata <= X"6BACA94D";
    when 16#17EB# => romdata <= X"37440049";
    when 16#17EC# => romdata <= X"9CA6813C";
    when 16#17ED# => romdata <= X"90A03DFE";
    when 16#17EE# => romdata <= X"2C537261";
    when 16#17EF# => romdata <= X"DA93A1C0";
    when 16#17F0# => romdata <= X"F6D8BA93";
    when 16#17F1# => romdata <= X"D1EB5FB1";
    when 16#17F2# => romdata <= X"7255DF28";
    when 16#17F3# => romdata <= X"B7873758";
    when 16#17F4# => romdata <= X"2FD675D0";
    when 16#17F5# => romdata <= X"56A4C474";
    when 16#17F6# => romdata <= X"A71CA8EF";
    when 16#17F7# => romdata <= X"0D77BAEB";
    when 16#17F8# => romdata <= X"E5637711";
    when 16#17F9# => romdata <= X"AEA3FF2B";
    when 16#17FA# => romdata <= X"01470044";
    when 16#17FB# => romdata <= X"8C3D74E3";
    when 16#17FC# => romdata <= X"DF264D77";
    when 16#17FD# => romdata <= X"3360F45C";
    when 16#17FE# => romdata <= X"CC334298";
    when 16#17FF# => romdata <= X"7169C9A0";
    when 16#1800# => romdata <= X"94741D7F";
    when 16#1801# => romdata <= X"05B0CA50";
    when 16#1802# => romdata <= X"908E6BC1";
    when 16#1803# => romdata <= X"4801A28E";
    when 16#1804# => romdata <= X"353551F0";
    when 16#1805# => romdata <= X"1769451B";
    when 16#1806# => romdata <= X"1482FAD0";
    when 16#1807# => romdata <= X"043D5C72";
    when 16#1808# => romdata <= X"331246D9";
    when 16#1809# => romdata <= X"AC3344F0";
    when 16#180A# => romdata <= X"FA2E28FD";
    when 16#180B# => romdata <= X"00E86B38";
    when 16#180C# => romdata <= X"F5E0452F";
    when 16#180D# => romdata <= X"46CA111E";
    when 16#180E# => romdata <= X"92D01B37";
    when 16#180F# => romdata <= X"E966455D";
    when 16#1810# => romdata <= X"F1374883";
    when 16#1811# => romdata <= X"DB8B055C";
    when 16#1812# => romdata <= X"4DF25B42";
    when 16#1813# => romdata <= X"182280F8";
    when 16#1814# => romdata <= X"6D0D825C";
    when 16#1815# => romdata <= X"096018D2";
    when 16#1816# => romdata <= X"949B4BFC";
    when 16#1817# => romdata <= X"EB7BB2C8";
    when 16#1818# => romdata <= X"A5BFA2C7";
    when 16#1819# => romdata <= X"9E27F11A";
    when 16#181A# => romdata <= X"7F9B43A5";
    when 16#181B# => romdata <= X"0AF928D8";
    when 16#181C# => romdata <= X"1FA95CEC";
    when 16#181D# => romdata <= X"86A11422";
    when 16#181E# => romdata <= X"2B997860";
    when 16#181F# => romdata <= X"72311025";
    when 16#1820# => romdata <= X"672AB04B";
    when 16#1821# => romdata <= X"2593C5AF";
    when 16#1822# => romdata <= X"50100B71";
    when 16#1823# => romdata <= X"D052AE26";
    when 16#1824# => romdata <= X"8FBA992B";
    when 16#1825# => romdata <= X"F7868E58";
    when 16#1826# => romdata <= X"EFCD07A2";
    when 16#1827# => romdata <= X"4D211177";
    when 16#1828# => romdata <= X"4A36115C";
    when 16#1829# => romdata <= X"1C527B51";
    when 16#182A# => romdata <= X"92EA9557";
    when 16#182B# => romdata <= X"22EAE849";
    when 16#182C# => romdata <= X"EF83817F";
    when 16#182D# => romdata <= X"E8595C96";
    when 16#182E# => romdata <= X"EA2D76FE";
    when 16#182F# => romdata <= X"CF6476D8";
    when 16#1830# => romdata <= X"9F65A262";
    when 16#1831# => romdata <= X"D94B3F5E";
    when 16#1832# => romdata <= X"89A5DE8B";
    when 16#1833# => romdata <= X"1A7333EF";
    when 16#1834# => romdata <= X"CDFDED17";
    when 16#1835# => romdata <= X"FE1CCADE";
    when 16#1836# => romdata <= X"BA0D1E7B";
    when 16#1837# => romdata <= X"73E67491";
    when 16#1838# => romdata <= X"B413A862";
    when 16#1839# => romdata <= X"E34A308D";
    when 16#183A# => romdata <= X"5C211787";
    when 16#183B# => romdata <= X"E6ED8683";
    when 16#183C# => romdata <= X"C6E1DDEB";
    when 16#183D# => romdata <= X"8EE2D281";
    when 16#183E# => romdata <= X"166C03E7";
    when 16#183F# => romdata <= X"A72D7D7B";
    when 16#1840# => romdata <= X"D8B878D0";
    when 16#1841# => romdata <= X"7D2216C2";
    when 16#1842# => romdata <= X"1B855CCD";
    when 16#1843# => romdata <= X"A76B7B75";
    when 16#1844# => romdata <= X"DD1B2CB8";
    when 16#1845# => romdata <= X"76E59F91";
    when 16#1846# => romdata <= X"F040D42B";
    when 16#1847# => romdata <= X"97050043";
    when 16#1848# => romdata <= X"499DCFFC";
    when 16#1849# => romdata <= X"65AF803E";
    when 16#184A# => romdata <= X"2F7455C9";
    when 16#184B# => romdata <= X"669DD989";
    when 16#184C# => romdata <= X"6FE1F622";
    when 16#184D# => romdata <= X"27936DF9";
    when 16#184E# => romdata <= X"05835A64";
    when 16#184F# => romdata <= X"4D31130A";
    when 16#1850# => romdata <= X"39479DE7";
    when 16#1851# => romdata <= X"5B4DC436";
    when 16#1852# => romdata <= X"1E41202D";
    when 16#1853# => romdata <= X"51D50E0E";
    when 16#1854# => romdata <= X"4B4B218A";
    when 16#1855# => romdata <= X"F7F5CAF2";
    when 16#1856# => romdata <= X"64DCD060";
    when 16#1857# => romdata <= X"C296E777";
    when 16#1858# => romdata <= X"DF1EED6A";
    when 16#1859# => romdata <= X"E8147E9B";
    when 16#185A# => romdata <= X"6CA73184";
    when 16#185B# => romdata <= X"C345FBDD";
    when 16#185C# => romdata <= X"89DE4A99";
    when 16#185D# => romdata <= X"9C42AB46";
    when 16#185E# => romdata <= X"81D9EA3B";
    when 16#185F# => romdata <= X"86DD7503";
    when 16#1860# => romdata <= X"1A33DCDC";
    when 16#1861# => romdata <= X"807F8FB1";
    when 16#1862# => romdata <= X"4EE0CE61";
    when 16#1863# => romdata <= X"B16068AF";
    when 16#1864# => romdata <= X"01CCE737";
    when 16#1865# => romdata <= X"8C9D9659";
    when 16#1866# => romdata <= X"43476AD2";
    when 16#1867# => romdata <= X"1A469D8B";
    when 16#1868# => romdata <= X"0CAE15BA";
    when 16#1869# => romdata <= X"8FE04971";
    when 16#186A# => romdata <= X"FE1EC61D";
    when 16#186B# => romdata <= X"3AAD3386";
    when 16#186C# => romdata <= X"DF71B33F";
    when 16#186D# => romdata <= X"D0B4F324";
    when 16#186E# => romdata <= X"F3DA518F";
    when 16#186F# => romdata <= X"0CC03531";
    when 16#1870# => romdata <= X"82B3D76C";
    when 16#1871# => romdata <= X"F4EF5AB1";
    when 16#1872# => romdata <= X"50FB9E74";
    when 16#1873# => romdata <= X"C28234CB";
    when 16#1874# => romdata <= X"3D907AC8";
    when 16#1875# => romdata <= X"1CB6D3B9";
    when 16#1876# => romdata <= X"9D510B48";
    when 16#1877# => romdata <= X"1E1F0423";
    when 16#1878# => romdata <= X"D6F4987F";
    when 16#1879# => romdata <= X"5517ABBB";
    when 16#187A# => romdata <= X"EEC07F46";
    when 16#187B# => romdata <= X"AECEBA5F";
    when 16#187C# => romdata <= X"15D91AEB";
    when 16#187D# => romdata <= X"0FE91490";
    when 16#187E# => romdata <= X"E91F739D";
    when 16#187F# => romdata <= X"465225C0";
    when 16#1880# => romdata <= X"839A0146";
    when 16#1881# => romdata <= X"4B473A64";
    when 16#1882# => romdata <= X"A3D1EA24";
    when 16#1883# => romdata <= X"EB363EAA";
    when 16#1884# => romdata <= X"A590F4BD";
    when 16#1885# => romdata <= X"0E4492FE";
    when 16#1886# => romdata <= X"C4E3D4DB";
    when 16#1887# => romdata <= X"5883E487";
    when 16#1888# => romdata <= X"3BBA1759";
    when 16#1889# => romdata <= X"5FF48134";
    when 16#188A# => romdata <= X"893F16F5";
    when 16#188B# => romdata <= X"C4A43659";
    when 16#188C# => romdata <= X"C46484A2";
    when 16#188D# => romdata <= X"68C3303B";
    when 16#188E# => romdata <= X"2DC345E8";
    when 16#188F# => romdata <= X"C98FBBA6";
    when 16#1890# => romdata <= X"D06946F9";
    when 16#1891# => romdata <= X"97074AE1";
    when 16#1892# => romdata <= X"5680EC94";
    when 16#1893# => romdata <= X"23D64645";
    when 16#1894# => romdata <= X"85D98804";
    when 16#1895# => romdata <= X"B3541662";
    when 16#1896# => romdata <= X"E183F654";
    when 16#1897# => romdata <= X"0503BEC2";
    when 16#1898# => romdata <= X"04749D58";
    when 16#1899# => romdata <= X"E3DB9ECF";
    when 16#189A# => romdata <= X"11C80CD3";
    when 16#189B# => romdata <= X"A38F8D66";
    when 16#189C# => romdata <= X"FFE6CC8A";
    when 16#189D# => romdata <= X"003BDD35";
    when 16#189E# => romdata <= X"F547E503";
    when 16#189F# => romdata <= X"9DE9A21F";
    when 16#18A0# => romdata <= X"70A8A07B";
    when 16#18A1# => romdata <= X"2DD89B68";
    when 16#18A2# => romdata <= X"E43B42C2";
    when 16#18A3# => romdata <= X"E021A119";
    when 16#18A4# => romdata <= X"09817C54";
    when 16#18A5# => romdata <= X"3F839E68";
    when 16#18A6# => romdata <= X"62268E38";
    when 16#18A7# => romdata <= X"DCE712B4";
    when 16#18A8# => romdata <= X"D49C39A5";
    when 16#18A9# => romdata <= X"035F3D6B";
    when 16#18AA# => romdata <= X"A19AE028";
    when 16#18AB# => romdata <= X"AE70CCF5";
    when 16#18AC# => romdata <= X"57720794";
    when 16#18AD# => romdata <= X"FEF64429";
    when 16#18AE# => romdata <= X"99E740CD";
    when 16#18AF# => romdata <= X"6AFE6235";
    when 16#18B0# => romdata <= X"F165515F";
    when 16#18B1# => romdata <= X"DC24AB6F";
    when 16#18B2# => romdata <= X"578DB254";
    when 16#18B3# => romdata <= X"9C8065E0";
    when 16#18B4# => romdata <= X"08577FCF";
    when 16#18B5# => romdata <= X"8B8DD8A3";
    when 16#18B6# => romdata <= X"BA679BAB";
    when 16#18B7# => romdata <= X"BC9A747A";
    when 16#18B8# => romdata <= X"4E2DABD9";
    when 16#18B9# => romdata <= X"1501424E";
    when 16#18BA# => romdata <= X"4191097E";
    when 16#18BB# => romdata <= X"689A741E";
    when 16#18BC# => romdata <= X"B6644A77";
    when 16#18BD# => romdata <= X"1CABDBFE";
    when 16#18BE# => romdata <= X"6B74ED3E";
    when 16#18BF# => romdata <= X"D171DF8D";
    when 16#18C0# => romdata <= X"E641C1D4";
    when 16#18C1# => romdata <= X"2213B9D0";
    when 16#18C2# => romdata <= X"F8CAD1E1";
    when 16#18C3# => romdata <= X"1FF63670";
    when 16#18C4# => romdata <= X"F5587F1F";
    when 16#18C5# => romdata <= X"B7FF9227";
    when 16#18C6# => romdata <= X"6AB48F31";
    when 16#18C7# => romdata <= X"751E7A59";
    when 16#18C8# => romdata <= X"1AF4F096";
    when 16#18C9# => romdata <= X"6F390988";
    when 16#18CA# => romdata <= X"3EE60156";
    when 16#18CB# => romdata <= X"39671BDC";
    when 16#18CC# => romdata <= X"3D137875";
    when 16#18CD# => romdata <= X"0F66F5DD";
    when 16#18CE# => romdata <= X"165912CF";
    when 16#18CF# => romdata <= X"F1A54ED4";
    when 16#18D0# => romdata <= X"63905404";
    when 16#18D1# => romdata <= X"EB7D3412";
    when 16#18D2# => romdata <= X"EE2B0F0D";
    when 16#18D3# => romdata <= X"9E6B99EC";
    when 16#18D4# => romdata <= X"81678ABC";
    when 16#18D5# => romdata <= X"D1789BD8";
    when 16#18D6# => romdata <= X"F1D72D3D";
    when 16#18D7# => romdata <= X"F8754A16";
    when 16#18D8# => romdata <= X"DC2106B8";
    when 16#18D9# => romdata <= X"3B325807";
    when 16#18DA# => romdata <= X"E27BCBD2";
    when 16#18DB# => romdata <= X"2A25DAC3";
    when 16#18DC# => romdata <= X"2F27EACA";
    when 16#18DD# => romdata <= X"B6A4CB6C";
    when 16#18DE# => romdata <= X"BA4CC90D";
    when 16#18DF# => romdata <= X"5302BE5E";
    when 16#18E0# => romdata <= X"9827B7AB";
    when 16#18E1# => romdata <= X"48BB696B";
    when 16#18E2# => romdata <= X"2902975C";
    when 16#18E3# => romdata <= X"48B3A4BA";
    when 16#18E4# => romdata <= X"4630B14E";
    when 16#18E5# => romdata <= X"0FD8A050";
    when 16#18E6# => romdata <= X"B0718C28";
    when 16#18E7# => romdata <= X"29371BEC";
    when 16#18E8# => romdata <= X"59738717";
    when 16#18E9# => romdata <= X"2B0B3192";
    when 16#18EA# => romdata <= X"EF958BD1";
    when 16#18EB# => romdata <= X"F7977EF9";
    when 16#18EC# => romdata <= X"A3A6C80D";
    when 16#18ED# => romdata <= X"53BC9613";
    when 16#18EE# => romdata <= X"15F97B71";
    when 16#18EF# => romdata <= X"4253B973";
    when 16#18F0# => romdata <= X"1A017BE2";
    when 16#18F1# => romdata <= X"CA1D4302";
    when 16#18F2# => romdata <= X"4F75E26B";
    when 16#18F3# => romdata <= X"BE989C4D";
    when 16#18F4# => romdata <= X"514D0153";
    when 16#18F5# => romdata <= X"8956FE4B";
    when 16#18F6# => romdata <= X"90BE17B3";
    when 16#18F7# => romdata <= X"407B55BD";
    when 16#18F8# => romdata <= X"08BA50FA";
    when 16#18F9# => romdata <= X"807D0E44";
    when 16#18FA# => romdata <= X"8B7CAC65";
    when 16#18FB# => romdata <= X"EB3FF856";
    when 16#18FC# => romdata <= X"772A933F";
    when 16#18FD# => romdata <= X"0C5F3E6F";
    when 16#18FE# => romdata <= X"41E05101";
    when 16#18FF# => romdata <= X"5C6F9B80";
    when 16#1900# => romdata <= X"BDA2B72F";
    when 16#1901# => romdata <= X"0BB02652";
    when 16#1902# => romdata <= X"69F19820";
    when 16#1903# => romdata <= X"7FB061DA";
    when 16#1904# => romdata <= X"29DE43E3";
    when 16#1905# => romdata <= X"0847E7C0";
    when 16#1906# => romdata <= X"62A581A7";
    when 16#1907# => romdata <= X"EB53491E";
    when 16#1908# => romdata <= X"A51B51ED";
    when 16#1909# => romdata <= X"D36F991D";
    when 16#190A# => romdata <= X"15AF89AB";
    when 16#190B# => romdata <= X"53198537";
    when 16#190C# => romdata <= X"988350FD";
    when 16#190D# => romdata <= X"5FDF8E00";
    when 16#190E# => romdata <= X"3019BE11";
    when 16#190F# => romdata <= X"5840B9BA";
    when 16#1910# => romdata <= X"55C238C3";
    when 16#1911# => romdata <= X"CBC72C0E";
    when 16#1912# => romdata <= X"24E25090";
    when 16#1913# => romdata <= X"A3D6A59B";
    when 16#1914# => romdata <= X"EA9FED0F";
    when 16#1915# => romdata <= X"AC9EAD40";
    when 16#1916# => romdata <= X"451A9564";
    when 16#1917# => romdata <= X"9638FE0B";
    when 16#1918# => romdata <= X"B0F8FFE6";
    when 16#1919# => romdata <= X"1AF5B9A8";
    when 16#191A# => romdata <= X"AB84BE84";
    when 16#191B# => romdata <= X"C65EA1E1";
    when 16#191C# => romdata <= X"2E9F6650";
    when 16#191D# => romdata <= X"ADB59A82";
    when 16#191E# => romdata <= X"4E608E80";
    when 16#191F# => romdata <= X"D1FC3AC1";
    when 16#1920# => romdata <= X"9F418169";
    when 16#1921# => romdata <= X"B3879CC9";
    when 16#1922# => romdata <= X"46165511";
    when 16#1923# => romdata <= X"D5AA280A";
    when 16#1924# => romdata <= X"E644AF36";
    when 16#1925# => romdata <= X"0C42F7A3";
    when 16#1926# => romdata <= X"EEDF27E3";
    when 16#1927# => romdata <= X"68E46480";
    when 16#1928# => romdata <= X"E3353E67";
    when 16#1929# => romdata <= X"F536E02B";
    when 16#192A# => romdata <= X"33505341";
    when 16#192B# => romdata <= X"BAF39410";
    when 16#192C# => romdata <= X"69567B72";
    when 16#192D# => romdata <= X"3D7C125C";
    when 16#192E# => romdata <= X"8F066F9A";
    when 16#192F# => romdata <= X"6255436A";
    when 16#1930# => romdata <= X"AFDCAA8C";
    when 16#1931# => romdata <= X"554FDAFB";
    when 16#1932# => romdata <= X"0A9AAD91";
    when 16#1933# => romdata <= X"F1263DC6";
    when 16#1934# => romdata <= X"2EF91A74";
    when 16#1935# => romdata <= X"8FFB29F5";
    when 16#1936# => romdata <= X"7E325D65";
    when 16#1937# => romdata <= X"A38ECB4F";
    when 16#1938# => romdata <= X"2851923D";
    when 16#1939# => romdata <= X"C6E9B729";
    when 16#193A# => romdata <= X"6064148A";
    when 16#193B# => romdata <= X"9BA2D938";
    when 16#193C# => romdata <= X"116266C5";
    when 16#193D# => romdata <= X"97D9E1F1";
    when 16#193E# => romdata <= X"1A46BE0E";
    when 16#193F# => romdata <= X"F526225B";
    when 16#1940# => romdata <= X"E750F0F3";
    when 16#1941# => romdata <= X"E5B0AEB7";
    when 16#1942# => romdata <= X"DC2140FA";
    when 16#1943# => romdata <= X"3A48B723";
    when 16#1944# => romdata <= X"8D0F5A87";
    when 16#1945# => romdata <= X"2000782C";
    when 16#1946# => romdata <= X"B6F77514";
    when 16#1947# => romdata <= X"43EC6A1B";
    when 16#1948# => romdata <= X"7FA1ED02";
    when 16#1949# => romdata <= X"B9ABCD1C";
    when 16#194A# => romdata <= X"1DE4FC85";
    when 16#194B# => romdata <= X"E9B405C7";
    when 16#194C# => romdata <= X"851913C6";
    when 16#194D# => romdata <= X"0F85582B";
    when 16#194E# => romdata <= X"1529276A";
    when 16#194F# => romdata <= X"D475AE52";
    when 16#1950# => romdata <= X"BD8115B6";
    when 16#1951# => romdata <= X"E73A5350";
    when 16#1952# => romdata <= X"6E7A0244";
    when 16#1953# => romdata <= X"E1C29BCE";
    when 16#1954# => romdata <= X"F4CF20CF";
    when 16#1955# => romdata <= X"DF883392";
    when 16#1956# => romdata <= X"BB3990BE";
    when 16#1957# => romdata <= X"2A11B321";
    when 16#1958# => romdata <= X"3B68EC4A";
    when 16#1959# => romdata <= X"166C77D7";
    when 16#195A# => romdata <= X"24CFAEBD";
    when 16#195B# => romdata <= X"C34C45ED";
    when 16#195C# => romdata <= X"09848A99";
    when 16#195D# => romdata <= X"4BCE1FF6";
    when 16#195E# => romdata <= X"A9BB80C7";
    when 16#195F# => romdata <= X"F5CA8FD4";
    when 16#1960# => romdata <= X"4D3FDF8D";
    when 16#1961# => romdata <= X"EC8BA655";
    when 16#1962# => romdata <= X"2C234EF8";
    when 16#1963# => romdata <= X"DC52382D";
    when 16#1964# => romdata <= X"52D2B01B";
    when 16#1965# => romdata <= X"B23404FC";
    when 16#1966# => romdata <= X"453725C7";
    when 16#1967# => romdata <= X"C9269A78";
    when 16#1968# => romdata <= X"5FE09C71";
    when 16#1969# => romdata <= X"2D4ADE70";
    when 16#196A# => romdata <= X"72B66295";
    when 16#196B# => romdata <= X"CA0C6405";
    when 16#196C# => romdata <= X"D9859E13";
    when 16#196D# => romdata <= X"4FBBD373";
    when 16#196E# => romdata <= X"7F2956DD";
    when 16#196F# => romdata <= X"1D718A9F";
    when 16#1970# => romdata <= X"8242CE95";
    when 16#1971# => romdata <= X"BDB1E49F";
    when 16#1972# => romdata <= X"265EBF19";
    when 16#1973# => romdata <= X"976BC46E";
    when 16#1974# => romdata <= X"29F7DE0E";
    when 16#1975# => romdata <= X"E5C89A43";
    when 16#1976# => romdata <= X"AF2E1075";
    when 16#1977# => romdata <= X"88A46E1B";
    when 16#1978# => romdata <= X"6762E6F8";
    when 16#1979# => romdata <= X"E48B8FC4";
    when 16#197A# => romdata <= X"F4FF93EC";
    when 16#197B# => romdata <= X"60938B8E";
    when 16#197C# => romdata <= X"5C371902";
    when 16#197D# => romdata <= X"2C750C43";
    when 16#197E# => romdata <= X"09FC62AD";
    when 16#197F# => romdata <= X"A4E90280";
    when 16#1980# => romdata <= X"D240216C";
    when 16#1981# => romdata <= X"5C4A7074";
    when 16#1982# => romdata <= X"2CAA03AE";
    when 16#1983# => romdata <= X"910E8859";
    when 16#1984# => romdata <= X"C92E5A90";
    when 16#1985# => romdata <= X"A352CB8B";
    when 16#1986# => romdata <= X"45847BAC";
    when 16#1987# => romdata <= X"7793E1F7";
    when 16#1988# => romdata <= X"5720D449";
    when 16#1989# => romdata <= X"19E896AD";
    when 16#198A# => romdata <= X"4581E1FD";
    when 16#198B# => romdata <= X"83986FF2";
    when 16#198C# => romdata <= X"35C9834B";
    when 16#198D# => romdata <= X"EECAA155";
    when 16#198E# => romdata <= X"6794BE49";
    when 16#198F# => romdata <= X"033E79D4";
    when 16#1990# => romdata <= X"CCDB4DC6";
    when 16#1991# => romdata <= X"7C5200E8";
    when 16#1992# => romdata <= X"B6A3EE89";
    when 16#1993# => romdata <= X"1E700B34";
    when 16#1994# => romdata <= X"8CBF092E";
    when 16#1995# => romdata <= X"4D3FA5E6";
    when 16#1996# => romdata <= X"48B620E3";
    when 16#1997# => romdata <= X"4E491D7B";
    when 16#1998# => romdata <= X"628A1FE7";
    when 16#1999# => romdata <= X"E2C45586";
    when 16#199A# => romdata <= X"B6577E50";
    when 16#199B# => romdata <= X"788687F0";
    when 16#199C# => romdata <= X"858C10F7";
    when 16#199D# => romdata <= X"8F371B25";
    when 16#199E# => romdata <= X"C712ED27";
    when 16#199F# => romdata <= X"60C3D605";
    when 16#19A0# => romdata <= X"D4ED4F05";
    when 16#19A1# => romdata <= X"2E8B66FC";
    when 16#19A2# => romdata <= X"308D3ADD";
    when 16#19A3# => romdata <= X"4A9B86F0";
    when 16#19A4# => romdata <= X"0CE4257E";
    when 16#19A5# => romdata <= X"ED085EAE";
    when 16#19A6# => romdata <= X"95FBB1E1";
    when 16#19A7# => romdata <= X"13FCB42C";
    when 16#19A8# => romdata <= X"E12BB607";
    when 16#19A9# => romdata <= X"6178A209";
    when 16#19AA# => romdata <= X"03C55DA5";
    when 16#19AB# => romdata <= X"70EF8A25";
    when 16#19AC# => romdata <= X"BA7AC8B7";
    when 16#19AD# => romdata <= X"E134B8D4";
    when 16#19AE# => romdata <= X"E35AB172";
    when 16#19AF# => romdata <= X"CA33CC97";
    when 16#19B0# => romdata <= X"294A5E7E";
    when 16#19B1# => romdata <= X"579B9361";
    when 16#19B2# => romdata <= X"B92B49B6";
    when 16#19B3# => romdata <= X"3BB19827";
    when 16#19B4# => romdata <= X"40015DFE";
    when 16#19B5# => romdata <= X"C1688298";
    when 16#19B6# => romdata <= X"9C917F50";
    when 16#19B7# => romdata <= X"D5FDD916";
    when 16#19B8# => romdata <= X"6FE1001F";
    when 16#19B9# => romdata <= X"3282D3C5";
    when 16#19BA# => romdata <= X"4A28AC7F";
    when 16#19BB# => romdata <= X"D773CCC0";
    when 16#19BC# => romdata <= X"634AF7CD";
    when 16#19BD# => romdata <= X"F225F941";
    when 16#19BE# => romdata <= X"07C169D2";
    when 16#19BF# => romdata <= X"F2BB757E";
    when 16#19C0# => romdata <= X"EB55933C";
    when 16#19C1# => romdata <= X"CE0FF116";
    when 16#19C2# => romdata <= X"D7FFBA99";
    when 16#19C3# => romdata <= X"2F9A075A";
    when 16#19C4# => romdata <= X"2439CCB3";
    when 16#19C5# => romdata <= X"69D5B5DE";
    when 16#19C6# => romdata <= X"460CADC9";
    when 16#19C7# => romdata <= X"F8C81D98";
    when 16#19C8# => romdata <= X"E71651AE";
    when 16#19C9# => romdata <= X"BFC2A918";
    when 16#19CA# => romdata <= X"C551082D";
    when 16#19CB# => romdata <= X"85F75675";
    when 16#19CC# => romdata <= X"CDC8CCA1";
    when 16#19CD# => romdata <= X"D3E486CF";
    when 16#19CE# => romdata <= X"FB3B025D";
    when 16#19CF# => romdata <= X"27C8D67C";
    when 16#19D0# => romdata <= X"451FDFCF";
    when 16#19D1# => romdata <= X"59C3BFA1";
    when 16#19D2# => romdata <= X"63EB7911";
    when 16#19D3# => romdata <= X"52390E94";
    when 16#19D4# => romdata <= X"88C604B9";
    when 16#19D5# => romdata <= X"B8116C32";
    when 16#19D6# => romdata <= X"9453A98F";
    when 16#19D7# => romdata <= X"7A104527";
    when 16#19D8# => romdata <= X"BC677411";
    when 16#19D9# => romdata <= X"034CC496";
    when 16#19DA# => romdata <= X"86108E56";
    when 16#19DB# => romdata <= X"9B7595E1";
    when 16#19DC# => romdata <= X"DDC85918";
    when 16#19DD# => romdata <= X"D90BBCB3";
    when 16#19DE# => romdata <= X"37855860";
    when 16#19DF# => romdata <= X"D6E4718C";
    when 16#19E0# => romdata <= X"0679DAB6";
    when 16#19E1# => romdata <= X"982D23FC";
    when 16#19E2# => romdata <= X"B6648E85";
    when 16#19E3# => romdata <= X"61F44BCF";
    when 16#19E4# => romdata <= X"9B052D8B";
    when 16#19E5# => romdata <= X"58384523";
    when 16#19E6# => romdata <= X"BC592C9B";
    when 16#19E7# => romdata <= X"7F824B96";
    when 16#19E8# => romdata <= X"AD1A39AE";
    when 16#19E9# => romdata <= X"BD2232D6";
    when 16#19EA# => romdata <= X"D34DC171";
    when 16#19EB# => romdata <= X"E8FBF933";
    when 16#19EC# => romdata <= X"900960F2";
    when 16#19ED# => romdata <= X"07B55597";
    when 16#19EE# => romdata <= X"759D23E1";
    when 16#19EF# => romdata <= X"E7945075";
    when 16#19F0# => romdata <= X"86114228";
    when 16#19F1# => romdata <= X"A2FC100C";
    when 16#19F2# => romdata <= X"C200D2B8";
    when 16#19F3# => romdata <= X"62DF3F26";
    when 16#19F4# => romdata <= X"E6D1C937";
    when 16#19F5# => romdata <= X"0373FE16";
    when 16#19F6# => romdata <= X"5C326D8C";
    when 16#19F7# => romdata <= X"29FD2F0B";
    when 16#19F8# => romdata <= X"3071AFD5";
    when 16#19F9# => romdata <= X"215781BF";
    when 16#19FA# => romdata <= X"B589F605";
    when 16#19FB# => romdata <= X"263FF065";
    when 16#19FC# => romdata <= X"B7A5CA3F";
    when 16#19FD# => romdata <= X"6AA9DE3F";
    when 16#19FE# => romdata <= X"D8BF5589";
    when 16#19FF# => romdata <= X"BDE35260";
    when 16#1A00# => romdata <= X"8E7752C5";
    when 16#1A01# => romdata <= X"2805DD0A";
    when 16#1A02# => romdata <= X"723D61F0";
    when 16#1A03# => romdata <= X"BBE0122D";
    when 16#1A04# => romdata <= X"F576A42B";
    when 16#1A05# => romdata <= X"5AFDF9F1";
    when 16#1A06# => romdata <= X"96A766C9";
    when 16#1A07# => romdata <= X"B3BFE296";
    when 16#1A08# => romdata <= X"DC16A892";
    when 16#1A09# => romdata <= X"FAECEEDD";
    when 16#1A0A# => romdata <= X"8256D2B1";
    when 16#1A0B# => romdata <= X"AE6BFE54";
    when 16#1A0C# => romdata <= X"37D4A269";
    when 16#1A0D# => romdata <= X"1803043B";
    when 16#1A0E# => romdata <= X"59862B30";
    when 16#1A0F# => romdata <= X"D68E4FF9";
    when 16#1A10# => romdata <= X"4A0700D7";
    when 16#1A11# => romdata <= X"35CFE967";
    when 16#1A12# => romdata <= X"299724DA";
    when 16#1A13# => romdata <= X"9D680200";
    when 16#1A14# => romdata <= X"C898EED1";
    when 16#1A15# => romdata <= X"C785E7B8";
    when 16#1A16# => romdata <= X"CEB14F1D";
    when 16#1A17# => romdata <= X"CDC73FC6";
    when 16#1A18# => romdata <= X"25F9678B";
    when 16#1A19# => romdata <= X"40760358";
    when 16#1A1A# => romdata <= X"7220C2FD";
    when 16#1A1B# => romdata <= X"FE0A47E8";
    when 16#1A1C# => romdata <= X"2ADF36C2";
    when 16#1A1D# => romdata <= X"6F942797";
    when 16#1A1E# => romdata <= X"D608BA6B";
    when 16#1A1F# => romdata <= X"38A3AD1A";
    when 16#1A20# => romdata <= X"967315E1";
    when 16#1A21# => romdata <= X"F2D665B2";
    when 16#1A22# => romdata <= X"7D51E350";
    when 16#1A23# => romdata <= X"F075531A";
    when 16#1A24# => romdata <= X"179DB2EE";
    when 16#1A25# => romdata <= X"D55547EA";
    when 16#1A26# => romdata <= X"61761CD2";
    when 16#1A27# => romdata <= X"B3962FCB";
    when 16#1A28# => romdata <= X"34727911";
    when 16#1A29# => romdata <= X"7D1C7A75";
    when 16#1A2A# => romdata <= X"74B49FFE";
    when 16#1A2B# => romdata <= X"0991AF57";
    when 16#1A2C# => romdata <= X"2A2B0C96";
    when 16#1A2D# => romdata <= X"2A8A7980";
    when 16#1A2E# => romdata <= X"0CFD524A";
    when 16#1A2F# => romdata <= X"AF9E6401";
    when 16#1A30# => romdata <= X"C4456960";
    when 16#1A31# => romdata <= X"0F41F044";
    when 16#1A32# => romdata <= X"22DB891D";
    when 16#1A33# => romdata <= X"25B9F714";
    when 16#1A34# => romdata <= X"713086BB";
    when 16#1A35# => romdata <= X"FD0FB268";
    when 16#1A36# => romdata <= X"E66A4FB1";
    when 16#1A37# => romdata <= X"0C0ABEEB";
    when 16#1A38# => romdata <= X"31D0FBFB";
    when 16#1A39# => romdata <= X"A20B0E4F";
    when 16#1A3A# => romdata <= X"FF404051";
    when 16#1A3B# => romdata <= X"596FC6F6";
    when 16#1A3C# => romdata <= X"C8093AD0";
    when 16#1A3D# => romdata <= X"1807FA52";
    when 16#1A3E# => romdata <= X"041CD330";
    when 16#1A3F# => romdata <= X"07B205D1";
    when 16#1A40# => romdata <= X"5D47AF73";
    when 16#1A41# => romdata <= X"3966411A";
    when 16#1A42# => romdata <= X"36F4C7B8";
    when 16#1A43# => romdata <= X"46D0BE04";
    when 16#1A44# => romdata <= X"9ADC21B8";
    when 16#1A45# => romdata <= X"9EA4CE0F";
    when 16#1A46# => romdata <= X"BA414C00";
    when 16#1A47# => romdata <= X"5E66F36F";
    when 16#1A48# => romdata <= X"ACF3C43B";
    when 16#1A49# => romdata <= X"474D47DA";
    when 16#1A4A# => romdata <= X"D78AC114";
    when 16#1A4B# => romdata <= X"D0171C03";
    when 16#1A4C# => romdata <= X"1DFBE4A1";
    when 16#1A4D# => romdata <= X"5FE1A226";
    when 16#1A4E# => romdata <= X"03CD79B6";
    when 16#1A4F# => romdata <= X"BB448B67";
    when 16#1A50# => romdata <= X"A4DEDC97";
    when 16#1A51# => romdata <= X"262F7B86";
    when 16#1A52# => romdata <= X"9C54F385";
    when 16#1A53# => romdata <= X"F3682C74";
    when 16#1A54# => romdata <= X"4ED5AD6C";
    when 16#1A55# => romdata <= X"0B6E1679";
    when 16#1A56# => romdata <= X"3920E6B4";
    when 16#1A57# => romdata <= X"5A024010";
    when 16#1A58# => romdata <= X"896D5FEC";
    when 16#1A59# => romdata <= X"FA111CC9";
    when 16#1A5A# => romdata <= X"F0C34E72";
    when 16#1A5B# => romdata <= X"8B32F2C4";
    when 16#1A5C# => romdata <= X"D45B8AA6";
    when 16#1A5D# => romdata <= X"9B621AB9";
    when 16#1A5E# => romdata <= X"AC3D9D79";
    when 16#1A5F# => romdata <= X"B38BF205";
    when 16#1A60# => romdata <= X"E8D0D19F";
    when 16#1A61# => romdata <= X"AC44A76B";
    when 16#1A62# => romdata <= X"9F564452";
    when 16#1A63# => romdata <= X"6E06858F";
    when 16#1A64# => romdata <= X"76B3EE2D";
    when 16#1A65# => romdata <= X"74AEB197";
    when 16#1A66# => romdata <= X"1D6B6E68";
    when 16#1A67# => romdata <= X"B8377339";
    when 16#1A68# => romdata <= X"9AC32203";
    when 16#1A69# => romdata <= X"164564B1";
    when 16#1A6A# => romdata <= X"02B26C37";
    when 16#1A6B# => romdata <= X"0A9FEC67";
    when 16#1A6C# => romdata <= X"3C285AE0";
    when 16#1A6D# => romdata <= X"D1D3DF23";
    when 16#1A6E# => romdata <= X"9D48B649";
    when 16#1A6F# => romdata <= X"2B89846E";
    when 16#1A70# => romdata <= X"BED4618A";
    when 16#1A71# => romdata <= X"EC940DC6";
    when 16#1A72# => romdata <= X"2AF4C3FF";
    when 16#1A73# => romdata <= X"0D56FC9F";
    when 16#1A74# => romdata <= X"BE23EE3B";
    when 16#1A75# => romdata <= X"0A4890BA";
    when 16#1A76# => romdata <= X"2665A88E";
    when 16#1A77# => romdata <= X"9F40C4B6";
    when 16#1A78# => romdata <= X"A770F963";
    when 16#1A79# => romdata <= X"0234ED10";
    when 16#1A7A# => romdata <= X"A3A7FF3C";
    when 16#1A7B# => romdata <= X"5BCCBA83";
    when 16#1A7C# => romdata <= X"6F3EDC8B";
    when 16#1A7D# => romdata <= X"821AB18D";
    when 16#1A7E# => romdata <= X"4B1D51D9";
    when 16#1A7F# => romdata <= X"962C3280";
    when 16#1A80# => romdata <= X"E682E9D8";
    when 16#1A81# => romdata <= X"E92A7837";
    when 16#1A82# => romdata <= X"823C9B77";
    when 16#1A83# => romdata <= X"14D267F9";
    when 16#1A84# => romdata <= X"CE290E9F";
    when 16#1A85# => romdata <= X"A6CC0A84";
    when 16#1A86# => romdata <= X"32D3F750";
    when 16#1A87# => romdata <= X"7DAF6CF6";
    when 16#1A88# => romdata <= X"81246AA4";
    when 16#1A89# => romdata <= X"C2323C6B";
    when 16#1A8A# => romdata <= X"53BCC6E5";
    when 16#1A8B# => romdata <= X"3B31F497";
    when 16#1A8C# => romdata <= X"42EE5F4E";
    when 16#1A8D# => romdata <= X"6F79DC36";
    when 16#1A8E# => romdata <= X"727E98B0";
    when 16#1A8F# => romdata <= X"6D0300ED";
    when 16#1A90# => romdata <= X"21F0CF5F";
    when 16#1A91# => romdata <= X"2B51D830";
    when 16#1A92# => romdata <= X"4A51D0B4";
    when 16#1A93# => romdata <= X"98F4BFA3";
    when 16#1A94# => romdata <= X"9C0049B8";
    when 16#1A95# => romdata <= X"117DAD33";
    when 16#1A96# => romdata <= X"4D4B2E37";
    when 16#1A97# => romdata <= X"676EC42D";
    when 16#1A98# => romdata <= X"FE0EED63";
    when 16#1A99# => romdata <= X"B3726872";
    when 16#1A9A# => romdata <= X"CCF9A102";
    when 16#1A9B# => romdata <= X"23A8A456";
    when 16#1A9C# => romdata <= X"3BE8AC26";
    when 16#1A9D# => romdata <= X"6E069700";
    when 16#1A9E# => romdata <= X"4921DCCE";
    when 16#1A9F# => romdata <= X"EA5DD80C";
    when 16#1AA0# => romdata <= X"62567FDE";
    when 16#1AA1# => romdata <= X"BF2AFDF0";
    when 16#1AA2# => romdata <= X"30192831";
    when 16#1AA3# => romdata <= X"A6FD871F";
    when 16#1AA4# => romdata <= X"63D5DADA";
    when 16#1AA5# => romdata <= X"4B270AA9";
    when 16#1AA6# => romdata <= X"EC0ACE47";
    when 16#1AA7# => romdata <= X"E75BD190";
    when 16#1AA8# => romdata <= X"18CB809B";
    when 16#1AA9# => romdata <= X"548D4F2C";
    when 16#1AAA# => romdata <= X"24831C38";
    when 16#1AAB# => romdata <= X"4DD2B807";
    when 16#1AAC# => romdata <= X"852F596B";
    when 16#1AAD# => romdata <= X"D4FE32CA";
    when 16#1AAE# => romdata <= X"B3A16899";
    when 16#1AAF# => romdata <= X"D0B100E9";
    when 16#1AB0# => romdata <= X"F96D06AA";
    when 16#1AB1# => romdata <= X"CB8DA8D5";
    when 16#1AB2# => romdata <= X"1DB0B0F6";
    when 16#1AB3# => romdata <= X"00F3B614";
    when 16#1AB4# => romdata <= X"461F5238";
    when 16#1AB5# => romdata <= X"188B5EDA";
    when 16#1AB6# => romdata <= X"68EA753B";
    when 16#1AB7# => romdata <= X"6ACC5856";
    when 16#1AB8# => romdata <= X"9E841BAF";
    when 16#1AB9# => romdata <= X"92CEE04E";
    when 16#1ABA# => romdata <= X"6E2626B1";
    when 16#1ABB# => romdata <= X"FBD01B9B";
    when 16#1ABC# => romdata <= X"67D1311B";
    when 16#1ABD# => romdata <= X"1C3D6742";
    when 16#1ABE# => romdata <= X"7298E2D1";
    when 16#1ABF# => romdata <= X"93F0647E";
    when 16#1AC0# => romdata <= X"A17D16FD";
    when 16#1AC1# => romdata <= X"7FD6A40A";
    when 16#1AC2# => romdata <= X"1BDBB320";
    when 16#1AC3# => romdata <= X"A1F5FC64";
    when 16#1AC4# => romdata <= X"B97759AF";
    when 16#1AC5# => romdata <= X"4EA92AAE";
    when 16#1AC6# => romdata <= X"B759B5DD";
    when 16#1AC7# => romdata <= X"30A726E9";
    when 16#1AC8# => romdata <= X"B8EAFA37";
    when 16#1AC9# => romdata <= X"2FBD83CB";
    when 16#1ACA# => romdata <= X"FF0000CA";
    when 16#1ACB# => romdata <= X"75F219A9";
    when 16#1ACC# => romdata <= X"5D6A3CDE";
    when 16#1ACD# => romdata <= X"38B8DFA9";
    when 16#1ACE# => romdata <= X"281609A2";
    when 16#1ACF# => romdata <= X"0EE39B73";
    when 16#1AD0# => romdata <= X"FEBDF6A1";
    when 16#1AD1# => romdata <= X"55359476";
    when 16#1AD2# => romdata <= X"D073E715";
    when 16#1AD3# => romdata <= X"3BC918C1";
    when 16#1AD4# => romdata <= X"191C9BAA";
    when 16#1AD5# => romdata <= X"F0E0F161";
    when 16#1AD6# => romdata <= X"384DAD8A";
    when 16#1AD7# => romdata <= X"FC31A3FC";
    when 16#1AD8# => romdata <= X"1E9EAFA4";
    when 16#1AD9# => romdata <= X"95E22D18";
    when 16#1ADA# => romdata <= X"C05194EB";
    when 16#1ADB# => romdata <= X"85298AB0";
    when 16#1ADC# => romdata <= X"F042E447";
    when 16#1ADD# => romdata <= X"DD627904";
    when 16#1ADE# => romdata <= X"B73E6E50";
    when 16#1ADF# => romdata <= X"5712DF01";
    when 16#1AE0# => romdata <= X"0531C88E";
    when 16#1AE1# => romdata <= X"695F6510";
    when 16#1AE2# => romdata <= X"C78B443C";
    when 16#1AE3# => romdata <= X"731D7FDC";
    when 16#1AE4# => romdata <= X"D62EB7C4";
    when 16#1AE5# => romdata <= X"015AB5D5";
    when 16#1AE6# => romdata <= X"30BD09CE";
    when 16#1AE7# => romdata <= X"5229FA4D";
    when 16#1AE8# => romdata <= X"C5642AF1";
    when 16#1AE9# => romdata <= X"76C39D60";
    when 16#1AEA# => romdata <= X"FE070DF6";
    when 16#1AEB# => romdata <= X"35CC5435";
    when 16#1AEC# => romdata <= X"136C7BB9";
    when 16#1AED# => romdata <= X"C4DC83B0";
    when 16#1AEE# => romdata <= X"D382B9BB";
    when 16#1AEF# => romdata <= X"636A6C2B";
    when 16#1AF0# => romdata <= X"38385429";
    when 16#1AF1# => romdata <= X"04D53B86";
    when 16#1AF2# => romdata <= X"2585FE6E";
    when 16#1AF3# => romdata <= X"C8960A9A";
    when 16#1AF4# => romdata <= X"77783D17";
    when 16#1AF5# => romdata <= X"B2D90506";
    when 16#1AF6# => romdata <= X"F5D60998";
    when 16#1AF7# => romdata <= X"602AE543";
    when 16#1AF8# => romdata <= X"0E86025C";
    when 16#1AF9# => romdata <= X"8864883C";
    when 16#1AFA# => romdata <= X"ECD7CE51";
    when 16#1AFB# => romdata <= X"B49CC295";
    when 16#1AFC# => romdata <= X"3A2A41D7";
    when 16#1AFD# => romdata <= X"EF8027F1";
    when 16#1AFE# => romdata <= X"A83815BB";
    when 16#1AFF# => romdata <= X"EF6F6B20";
    when 16#1B00# => romdata <= X"F6BD4204";
    when 16#1B01# => romdata <= X"243CBA14";
    when 16#1B02# => romdata <= X"DAA15A25";
    when 16#1B03# => romdata <= X"6FBCD138";
    when 16#1B04# => romdata <= X"B5D875E2";
    when 16#1B05# => romdata <= X"8BCC0BA3";
    when 16#1B06# => romdata <= X"6855E648";
    when 16#1B07# => romdata <= X"434CD04F";
    when 16#1B08# => romdata <= X"49935C3D";
    when 16#1B09# => romdata <= X"074DD5BA";
    when 16#1B0A# => romdata <= X"2EB82AB1";
    when 16#1B0B# => romdata <= X"4E82C309";
    when 16#1B0C# => romdata <= X"91A1159E";
    when 16#1B0D# => romdata <= X"990D1D36";
    when 16#1B0E# => romdata <= X"DAF79485";
    when 16#1B0F# => romdata <= X"3A23C499";
    when 16#1B10# => romdata <= X"AB6B3DC0";
    when 16#1B11# => romdata <= X"2A89F014";
    when 16#1B12# => romdata <= X"31037281";
    when 16#1B13# => romdata <= X"3643F786";
    when 16#1B14# => romdata <= X"BF19D3FA";
    when 16#1B15# => romdata <= X"8C463EE5";
    when 16#1B16# => romdata <= X"0D9FA871";
    when 16#1B17# => romdata <= X"07E91C46";
    when 16#1B18# => romdata <= X"1AD2E5DF";
    when 16#1B19# => romdata <= X"2FC99630";
    when 16#1B1A# => romdata <= X"D2005894";
    when 16#1B1B# => romdata <= X"CB769812";
    when 16#1B1C# => romdata <= X"3111FAFC";
    when 16#1B1D# => romdata <= X"0C5BC9D1";
    when 16#1B1E# => romdata <= X"E8E84FCC";
    when 16#1B1F# => romdata <= X"A5179A6C";
    when 16#1B20# => romdata <= X"9AFE3E36";
    when 16#1B21# => romdata <= X"9222D668";
    when 16#1B22# => romdata <= X"54F90D26";
    when 16#1B23# => romdata <= X"68A57FDE";
    when 16#1B24# => romdata <= X"E00C300A";
    when 16#1B25# => romdata <= X"EA4E88F0";
    when 16#1B26# => romdata <= X"3F05C4D7";
    when 16#1B27# => romdata <= X"695B206D";
    when 16#1B28# => romdata <= X"E9F7E1D4";
    when 16#1B29# => romdata <= X"29E5E6B6";
    when 16#1B2A# => romdata <= X"5DFE05D4";
    when 16#1B2B# => romdata <= X"C861F4E7";
    when 16#1B2C# => romdata <= X"844DDB90";
    when 16#1B2D# => romdata <= X"62C0B6DB";
    when 16#1B2E# => romdata <= X"46B27AD0";
    when 16#1B2F# => romdata <= X"368992F5";
    when 16#1B30# => romdata <= X"4A44829D";
    when 16#1B31# => romdata <= X"D11A05AB";
    when 16#1B32# => romdata <= X"97BA8AD8";
    when 16#1B33# => romdata <= X"54E428B8";
    when 16#1B34# => romdata <= X"7F20C4E5";
    when 16#1B35# => romdata <= X"E4BB1FF3";
    when 16#1B36# => romdata <= X"803809A8";
    when 16#1B37# => romdata <= X"1F2E4C10";
    when 16#1B38# => romdata <= X"95720067";
    when 16#1B39# => romdata <= X"29A5E490";
    when 16#1B3A# => romdata <= X"E0AA40BA";
    when 16#1B3B# => romdata <= X"55F4391C";
    when 16#1B3C# => romdata <= X"9FB758EF";
    when 16#1B3D# => romdata <= X"A79B97E6";
    when 16#1B3E# => romdata <= X"D413BCB0";
    when 16#1B3F# => romdata <= X"2D33A00D";
    when 16#1B40# => romdata <= X"A6705BFB";
    when 16#1B41# => romdata <= X"ADED66CF";
    when 16#1B42# => romdata <= X"C21291C4";
    when 16#1B43# => romdata <= X"94B7C329";
    when 16#1B44# => romdata <= X"3810012E";
    when 16#1B45# => romdata <= X"CC61415E";
    when 16#1B46# => romdata <= X"609DD97A";
    when 16#1B47# => romdata <= X"AFFDEB79";
    when 16#1B48# => romdata <= X"5DE36026";
    when 16#1B49# => romdata <= X"B4602DD5";
    when 16#1B4A# => romdata <= X"46A1AD93";
    when 16#1B4B# => romdata <= X"7F1A6DEA";
    when 16#1B4C# => romdata <= X"CD3393F5";
    when 16#1B4D# => romdata <= X"530C48A7";
    when 16#1B4E# => romdata <= X"974E2882";
    when 16#1B4F# => romdata <= X"CB327AE6";
    when 16#1B50# => romdata <= X"00C05A53";
    when 16#1B51# => romdata <= X"5BDE5D15";
    when 16#1B52# => romdata <= X"AC524859";
    when 16#1B53# => romdata <= X"582EEE2D";
    when 16#1B54# => romdata <= X"62194B73";
    when 16#1B55# => romdata <= X"E0164335";
    when 16#1B56# => romdata <= X"9E7B2625";
    when 16#1B57# => romdata <= X"F3EB9FE7";
    when 16#1B58# => romdata <= X"137514ED";
    when 16#1B59# => romdata <= X"549A3196";
    when 16#1B5A# => romdata <= X"FFCBC807";
    when 16#1B5B# => romdata <= X"2B4F6C18";
    when 16#1B5C# => romdata <= X"CC67AAFA";
    when 16#1B5D# => romdata <= X"0ED6029A";
    when 16#1B5E# => romdata <= X"805EF098";
    when 16#1B5F# => romdata <= X"7E2F27A3";
    when 16#1B60# => romdata <= X"260F849C";
    when 16#1B61# => romdata <= X"68F3EF91";
    when 16#1B62# => romdata <= X"DAA9E579";
    when 16#1B63# => romdata <= X"AA16FDA6";
    when 16#1B64# => romdata <= X"98CC18AE";
    when 16#1B65# => romdata <= X"8706E28C";
    when 16#1B66# => romdata <= X"6D84CB3F";
    when 16#1B67# => romdata <= X"593273D7";
    when 16#1B68# => romdata <= X"63C29699";
    when 16#1B69# => romdata <= X"33D8EFA5";
    when 16#1B6A# => romdata <= X"64E8C06C";
    when 16#1B6B# => romdata <= X"427809E6";
    when 16#1B6C# => romdata <= X"A5A6F76D";
    when 16#1B6D# => romdata <= X"E7C8B07F";
    when 16#1B6E# => romdata <= X"F4EDDF6C";
    when 16#1B6F# => romdata <= X"F2B75950";
    when 16#1B70# => romdata <= X"66DFB15F";
    when 16#1B71# => romdata <= X"5C6F3839";
    when 16#1B72# => romdata <= X"DEE642FC";
    when 16#1B73# => romdata <= X"86BC1F3A";
    when 16#1B74# => romdata <= X"ED7ED2E6";
    when 16#1B75# => romdata <= X"5B665198";
    when 16#1B76# => romdata <= X"AA034817";
    when 16#1B77# => romdata <= X"DBBBE0FE";
    when 16#1B78# => romdata <= X"30E662B2";
    when 16#1B79# => romdata <= X"161276CB";
    when 16#1B7A# => romdata <= X"D969FDA0";
    when 16#1B7B# => romdata <= X"5AFD6D6A";
    when 16#1B7C# => romdata <= X"570C1E3C";
    when 16#1B7D# => romdata <= X"F7E32463";
    when 16#1B7E# => romdata <= X"4441983F";
    when 16#1B7F# => romdata <= X"257E2BA0";
    when 16#1B80# => romdata <= X"A9366308";
    when 16#1B81# => romdata <= X"475F2D8D";
    when 16#1B82# => romdata <= X"0C2D451C";
    when 16#1B83# => romdata <= X"4A65A01E";
    when 16#1B84# => romdata <= X"E58A0AF1";
    when 16#1B85# => romdata <= X"9B791D97";
    when 16#1B86# => romdata <= X"382EC59A";
    when 16#1B87# => romdata <= X"52616C74";
    when 16#1B88# => romdata <= X"80B86EB1";
    when 16#1B89# => romdata <= X"D0A83E93";
    when 16#1B8A# => romdata <= X"224B0DF7";
    when 16#1B8B# => romdata <= X"3DE1D7EE";
    when 16#1B8C# => romdata <= X"6D51088F";
    when 16#1B8D# => romdata <= X"3B20B793";
    when 16#1B8E# => romdata <= X"7E6C0144";
    when 16#1B8F# => romdata <= X"E0DACA63";
    when 16#1B90# => romdata <= X"24F0C8E5";
    when 16#1B91# => romdata <= X"F9D93A8C";
    when 16#1B92# => romdata <= X"BA1045E5";
    when 16#1B93# => romdata <= X"B509D7DF";
    when 16#1B94# => romdata <= X"98619FDD";
    when 16#1B95# => romdata <= X"FDD7892C";
    when 16#1B96# => romdata <= X"3082D690";
    when 16#1B97# => romdata <= X"08D9D3ED";
    when 16#1B98# => romdata <= X"6C9C1367";
    when 16#1B99# => romdata <= X"D9DB7C04";
    when 16#1B9A# => romdata <= X"621D7CDD";
    when 16#1B9B# => romdata <= X"8A5A2599";
    when 16#1B9C# => romdata <= X"EE45B87A";
    when 16#1B9D# => romdata <= X"82F8CE8D";
    when 16#1B9E# => romdata <= X"60293E7A";
    when 16#1B9F# => romdata <= X"71D11700";
    when 16#1BA0# => romdata <= X"CA9AF117";
    when 16#1BA1# => romdata <= X"D630C5D8";
    when 16#1BA2# => romdata <= X"B876A9DC";
    when 16#1BA3# => romdata <= X"E519BD65";
    when 16#1BA4# => romdata <= X"3114448C";
    when 16#1BA5# => romdata <= X"68B26581";
    when 16#1BA6# => romdata <= X"3C608435";
    when 16#1BA7# => romdata <= X"B96CD642";
    when 16#1BA8# => romdata <= X"A420A15F";
    when 16#1BA9# => romdata <= X"BAB46769";
    when 16#1BAA# => romdata <= X"2931BCA7";
    when 16#1BAB# => romdata <= X"4F1F9D23";
    when 16#1BAC# => romdata <= X"F5BFDDC5";
    when 16#1BAD# => romdata <= X"B8651139";
    when 16#1BAE# => romdata <= X"B5A73F04";
    when 16#1BAF# => romdata <= X"FEF3DA64";
    when 16#1BB0# => romdata <= X"B7BD56E4";
    when 16#1BB1# => romdata <= X"9235069E";
    when 16#1BB2# => romdata <= X"E5E8A136";
    when 16#1BB3# => romdata <= X"B921051F";
    when 16#1BB4# => romdata <= X"1D1C7D59";
    when 16#1BB5# => romdata <= X"93E6EEEE";
    when 16#1BB6# => romdata <= X"A2D58583";
    when 16#1BB7# => romdata <= X"152ADCD8";
    when 16#1BB8# => romdata <= X"7AA89CF5";
    when 16#1BB9# => romdata <= X"962BC834";
    when 16#1BBA# => romdata <= X"1EF99CEB";
    when 16#1BBB# => romdata <= X"3682A2D0";
    when 16#1BBC# => romdata <= X"686602CE";
    when 16#1BBD# => romdata <= X"140ABC2F";
    when 16#1BBE# => romdata <= X"DF79A778";
    when 16#1BBF# => romdata <= X"A9D75AFF";
    when 16#1BC0# => romdata <= X"DBBA00C0";
    when 16#1BC1# => romdata <= X"BD6A8A8A";
    when 16#1BC2# => romdata <= X"FF9B5D1F";
    when 16#1BC3# => romdata <= X"30C83735";
    when 16#1BC4# => romdata <= X"72C81BD9";
    when 16#1BC5# => romdata <= X"59489010";
    when 16#1BC6# => romdata <= X"2F46B5A3";
    when 16#1BC7# => romdata <= X"93ED126C";
    when 16#1BC8# => romdata <= X"36AEF6A6";
    when 16#1BC9# => romdata <= X"6E231A24";
    when 16#1BCA# => romdata <= X"6FDFCBD3";
    when 16#1BCB# => romdata <= X"DED198AB";
    when 16#1BCC# => romdata <= X"C54CF357";
    when 16#1BCD# => romdata <= X"ABC67AC8";
    when 16#1BCE# => romdata <= X"3680C048";
    when 16#1BCF# => romdata <= X"932D7C90";
    when 16#1BD0# => romdata <= X"2AB7DB16";
    when 16#1BD1# => romdata <= X"952B3C95";
    when 16#1BD2# => romdata <= X"DF4E845B";
    when 16#1BD3# => romdata <= X"46A362FF";
    when 16#1BD4# => romdata <= X"E1A27CD1";
    when 16#1BD5# => romdata <= X"388483FF";
    when 16#1BD6# => romdata <= X"A41AA563";
    when 16#1BD7# => romdata <= X"933371C0";
    when 16#1BD8# => romdata <= X"180848F9";
    when 16#1BD9# => romdata <= X"E3C03AFC";
    when 16#1BDA# => romdata <= X"1F00D6AB";
    when 16#1BDB# => romdata <= X"A29A9533";
    when 16#1BDC# => romdata <= X"27A4E3D9";
    when 16#1BDD# => romdata <= X"FAD4616C";
    when 16#1BDE# => romdata <= X"8546C9AF";
    when 16#1BDF# => romdata <= X"89FB4D08";
    when 16#1BE0# => romdata <= X"D4256923";
    when 16#1BE1# => romdata <= X"B736A8F6";
    when 16#1BE2# => romdata <= X"8FEA5A09";
    when 16#1BE3# => romdata <= X"7E0640C1";
    when 16#1BE4# => romdata <= X"6E0F7F94";
    when 16#1BE5# => romdata <= X"2E6A6F5C";
    when 16#1BE6# => romdata <= X"BA76BB00";
    when 16#1BE7# => romdata <= X"D81C606C";
    when 16#1BE8# => romdata <= X"7FED9087";
    when 16#1BE9# => romdata <= X"89A63F01";
    when 16#1BEA# => romdata <= X"F9B5FC7B";
    when 16#1BEB# => romdata <= X"7BE434E8";
    when 16#1BEC# => romdata <= X"5A0A44B2";
    when 16#1BED# => romdata <= X"070BE71A";
    when 16#1BEE# => romdata <= X"B2BA0132";
    when 16#1BEF# => romdata <= X"D9D7B32E";
    when 16#1BF0# => romdata <= X"2D2FE229";
    when 16#1BF1# => romdata <= X"619F8564";
    when 16#1BF2# => romdata <= X"3E75B414";
    when 16#1BF3# => romdata <= X"1D355386";
    when 16#1BF4# => romdata <= X"D1A09F45";
    when 16#1BF5# => romdata <= X"738455BC";
    when 16#1BF6# => romdata <= X"21607086";
    when 16#1BF7# => romdata <= X"C7BBCD4B";
    when 16#1BF8# => romdata <= X"73F87DD8";
    when 16#1BF9# => romdata <= X"3E905BCE";
    when 16#1BFA# => romdata <= X"8FC6C5BF";
    when 16#1BFB# => romdata <= X"1824E904";
    when 16#1BFC# => romdata <= X"C4F5C265";
    when 16#1BFD# => romdata <= X"18B2FEBF";
    when 16#1BFE# => romdata <= X"8EB06B22";
    when 16#1BFF# => romdata <= X"437270C0";
    when 16#1C00# => romdata <= X"92D87BF3";
    when 16#1C01# => romdata <= X"F54B0445";
    when 16#1C02# => romdata <= X"C05E508E";
    when 16#1C03# => romdata <= X"80F9CBC0";
    when 16#1C04# => romdata <= X"502F0897";
    when 16#1C05# => romdata <= X"D717CA23";
    when 16#1C06# => romdata <= X"2004362F";
    when 16#1C07# => romdata <= X"394A023B";
    when 16#1C08# => romdata <= X"FBFE3322";
    when 16#1C09# => romdata <= X"C1D331AF";
    when 16#1C0A# => romdata <= X"C6454FC7";
    when 16#1C0B# => romdata <= X"56FB4876";
    when 16#1C0C# => romdata <= X"8693FD5C";
    when 16#1C0D# => romdata <= X"46DDB40D";
    when 16#1C0E# => romdata <= X"CBF14C72";
    when 16#1C0F# => romdata <= X"6C24ED67";
    when 16#1C10# => romdata <= X"D8F3EB61";
    when 16#1C11# => romdata <= X"3BA80B0E";
    when 16#1C12# => romdata <= X"39CF0747";
    when 16#1C13# => romdata <= X"DF62D258";
    when 16#1C14# => romdata <= X"613640D8";
    when 16#1C15# => romdata <= X"81E085C3";
    when 16#1C16# => romdata <= X"77DE1C3D";
    when 16#1C17# => romdata <= X"149C8359";
    when 16#1C18# => romdata <= X"407C2C6A";
    when 16#1C19# => romdata <= X"BC0D2718";
    when 16#1C1A# => romdata <= X"A2D42439";
    when 16#1C1B# => romdata <= X"A8E7B38C";
    when 16#1C1C# => romdata <= X"D7DCED72";
    when 16#1C1D# => romdata <= X"AE750B2B";
    when 16#1C1E# => romdata <= X"E88D0069";
    when 16#1C1F# => romdata <= X"FBE94BD6";
    when 16#1C20# => romdata <= X"9A9A4B4A";
    when 16#1C21# => romdata <= X"D42FEC5E";
    when 16#1C22# => romdata <= X"651A31F8";
    when 16#1C23# => romdata <= X"6B90DC2F";
    when 16#1C24# => romdata <= X"EBAA6FA6";
    when 16#1C25# => romdata <= X"E5F6368B";
    when 16#1C26# => romdata <= X"620C1750";
    when 16#1C27# => romdata <= X"278DF393";
    when 16#1C28# => romdata <= X"F7C5035D";
    when 16#1C29# => romdata <= X"47897FC0";
    when 16#1C2A# => romdata <= X"5FBC419A";
    when 16#1C2B# => romdata <= X"61330135";
    when 16#1C2C# => romdata <= X"F24365F1";
    when 16#1C2D# => romdata <= X"3D653D77";
    when 16#1C2E# => romdata <= X"CA2930DB";
    when 16#1C2F# => romdata <= X"B05A3815";
    when 16#1C30# => romdata <= X"FE83F75B";
    when 16#1C31# => romdata <= X"B1BD8B2D";
    when 16#1C32# => romdata <= X"E12A2FAA";
    when 16#1C33# => romdata <= X"DCD1ED62";
    when 16#1C34# => romdata <= X"329C55B8";
    when 16#1C35# => romdata <= X"7FB32CC8";
    when 16#1C36# => romdata <= X"F3B42D88";
    when 16#1C37# => romdata <= X"8981B419";
    when 16#1C38# => romdata <= X"2480D1F5";
    when 16#1C39# => romdata <= X"7CEB0C55";
    when 16#1C3A# => romdata <= X"897BDA6B";
    when 16#1C3B# => romdata <= X"9C0ACE1E";
    when 16#1C3C# => romdata <= X"7E4595E3";
    when 16#1C3D# => romdata <= X"0C736830";
    when 16#1C3E# => romdata <= X"62432084";
    when 16#1C3F# => romdata <= X"44FCF457";
    when 16#1C40# => romdata <= X"4C47B077";
    when 16#1C41# => romdata <= X"25B25EC2";
    when 16#1C42# => romdata <= X"E28F4C50";
    when 16#1C43# => romdata <= X"B744B386";
    when 16#1C44# => romdata <= X"0B361DDD";
    when 16#1C45# => romdata <= X"D22D949A";
    when 16#1C46# => romdata <= X"A94EBA4F";
    when 16#1C47# => romdata <= X"97606FCA";
    when 16#1C48# => romdata <= X"D91394B6";
    when 16#1C49# => romdata <= X"FC0E634B";
    when 16#1C4A# => romdata <= X"D15E099E";
    when 16#1C4B# => romdata <= X"697403B2";
    when 16#1C4C# => romdata <= X"AE84CDF5";
    when 16#1C4D# => romdata <= X"DBDF36D9";
    when 16#1C4E# => romdata <= X"1FB82C0B";
    when 16#1C4F# => romdata <= X"C12B984F";
    when 16#1C50# => romdata <= X"EE83CA9E";
    when 16#1C51# => romdata <= X"97C194CA";
    when 16#1C52# => romdata <= X"DF8382CE";
    when 16#1C53# => romdata <= X"CAAF49EB";
    when 16#1C54# => romdata <= X"3BD446F6";
    when 16#1C55# => romdata <= X"60F94C18";
    when 16#1C56# => romdata <= X"8C074CC3";
    when 16#1C57# => romdata <= X"12E186BE";
    when 16#1C58# => romdata <= X"E0F65855";
    when 16#1C59# => romdata <= X"35B050C2";
    when 16#1C5A# => romdata <= X"26659A94";
    when 16#1C5B# => romdata <= X"B4C4974D";
    when 16#1C5C# => romdata <= X"A32CDFF3";
    when 16#1C5D# => romdata <= X"0DBEB4DE";
    when 16#1C5E# => romdata <= X"A588C6F4";
    when 16#1C5F# => romdata <= X"90F7432D";
    when 16#1C60# => romdata <= X"A5FA2408";
    when 16#1C61# => romdata <= X"BBC931EA";
    when 16#1C62# => romdata <= X"F60EADD7";
    when 16#1C63# => romdata <= X"B891A61C";
    when 16#1C64# => romdata <= X"157147B8";
    when 16#1C65# => romdata <= X"DDE7A45F";
    when 16#1C66# => romdata <= X"909BD20D";
    when 16#1C67# => romdata <= X"5B120097";
    when 16#1C68# => romdata <= X"83DE4109";
    when 16#1C69# => romdata <= X"40245FE4";
    when 16#1C6A# => romdata <= X"E91ACCF7";
    when 16#1C6B# => romdata <= X"2942E486";
    when 16#1C6C# => romdata <= X"AE773CD6";
    when 16#1C6D# => romdata <= X"65912173";
    when 16#1C6E# => romdata <= X"EA29875A";
    when 16#1C6F# => romdata <= X"1722F865";
    when 16#1C70# => romdata <= X"8C414CD0";
    when 16#1C71# => romdata <= X"8CBFDFE1";
    when 16#1C72# => romdata <= X"DD356E16";
    when 16#1C73# => romdata <= X"7A9D7B20";
    when 16#1C74# => romdata <= X"BF744156";
    when 16#1C75# => romdata <= X"2EE81643";
    when 16#1C76# => romdata <= X"5A78BAE7";
    when 16#1C77# => romdata <= X"E5A5EB4D";
    when 16#1C78# => romdata <= X"A6AAAC36";
    when 16#1C79# => romdata <= X"F594C93E";
    when 16#1C7A# => romdata <= X"2851D76B";
    when 16#1C7B# => romdata <= X"6A18B0B0";
    when 16#1C7C# => romdata <= X"3B30CD38";
    when 16#1C7D# => romdata <= X"B97E3810";
    when 16#1C7E# => romdata <= X"9C494C55";
    when 16#1C7F# => romdata <= X"7643D580";
    when 16#1C80# => romdata <= X"BAA2716F";
    when 16#1C81# => romdata <= X"115D72D2";
    when 16#1C82# => romdata <= X"037841EF";
    when 16#1C83# => romdata <= X"9138D198";
    when 16#1C84# => romdata <= X"33C7C5FF";
    when 16#1C85# => romdata <= X"40F058A9";
    when 16#1C86# => romdata <= X"60826E69";
    when 16#1C87# => romdata <= X"03155777";
    when 16#1C88# => romdata <= X"10EFE64B";
    when 16#1C89# => romdata <= X"B3769156";
    when 16#1C8A# => romdata <= X"4B3B0B6C";
    when 16#1C8B# => romdata <= X"577DA603";
    when 16#1C8C# => romdata <= X"CC3ACDFE";
    when 16#1C8D# => romdata <= X"1785541A";
    when 16#1C8E# => romdata <= X"AD239047";
    when 16#1C8F# => romdata <= X"58A5A13B";
    when 16#1C90# => romdata <= X"DB018E71";
    when 16#1C91# => romdata <= X"69D479A1";
    when 16#1C92# => romdata <= X"FAA031CA";
    when 16#1C93# => romdata <= X"72FA6D6A";
    when 16#1C94# => romdata <= X"E9613D6B";
    when 16#1C95# => romdata <= X"2F82AB07";
    when 16#1C96# => romdata <= X"500B49DF";
    when 16#1C97# => romdata <= X"535F86A7";
    when 16#1C98# => romdata <= X"6350C140";
    when 16#1C99# => romdata <= X"F9CD2529";
    when 16#1C9A# => romdata <= X"5D6BC2F3";
    when 16#1C9B# => romdata <= X"8C5D13C9";
    when 16#1C9C# => romdata <= X"9540E236";
    when 16#1C9D# => romdata <= X"3862F06D";
    when 16#1C9E# => romdata <= X"DCC486D8";
    when 16#1C9F# => romdata <= X"84999BCB";
    when 16#1CA0# => romdata <= X"840BCCAF";
    when 16#1CA1# => romdata <= X"2AB84F59";
    when 16#1CA2# => romdata <= X"06B9AA0F";
    when 16#1CA3# => romdata <= X"77D6432F";
    when 16#1CA4# => romdata <= X"65315583";
    when 16#1CA5# => romdata <= X"92641C52";
    when 16#1CA6# => romdata <= X"FEAF9D8E";
    when 16#1CA7# => romdata <= X"D86BF015";
    when 16#1CA8# => romdata <= X"8134129F";
    when 16#1CA9# => romdata <= X"34ECD076";
    when 16#1CAA# => romdata <= X"8BC02ED4";
    when 16#1CAB# => romdata <= X"42254515";
    when 16#1CAC# => romdata <= X"A74999C6";
    when 16#1CAD# => romdata <= X"B8052A1F";
    when 16#1CAE# => romdata <= X"C797F572";
    when 16#1CAF# => romdata <= X"0738C69D";
    when 16#1CB0# => romdata <= X"D9B3FFAB";
    when 16#1CB1# => romdata <= X"DDC8515C";
    when 16#1CB2# => romdata <= X"D279B246";
    when 16#1CB3# => romdata <= X"EA7C6775";
    when 16#1CB4# => romdata <= X"4920038C";
    when 16#1CB5# => romdata <= X"5A4C8D30";
    when 16#1CB6# => romdata <= X"1119CEB9";
    when 16#1CB7# => romdata <= X"5FAB2765";
    when 16#1CB8# => romdata <= X"DE39DDA8";
    when 16#1CB9# => romdata <= X"4180CEBA";
    when 16#1CBA# => romdata <= X"AFBF4976";
    when 16#1CBB# => romdata <= X"118A8373";
    when 16#1CBC# => romdata <= X"FF6BBFC7";
    when 16#1CBD# => romdata <= X"FEBC3CFE";
    when 16#1CBE# => romdata <= X"AB1DA69D";
    when 16#1CBF# => romdata <= X"D3DB9E42";
    when 16#1CC0# => romdata <= X"8C594950";
    when 16#1CC1# => romdata <= X"FD51F4D9";
    when 16#1CC2# => romdata <= X"8A393BAB";
    when 16#1CC3# => romdata <= X"96001461";
    when 16#1CC4# => romdata <= X"F2765834";
    when 16#1CC5# => romdata <= X"ED70C60B";
    when 16#1CC6# => romdata <= X"C56406CF";
    when 16#1CC7# => romdata <= X"CB3E784C";
    when 16#1CC8# => romdata <= X"59B91C19";
    when 16#1CC9# => romdata <= X"783E67CE";
    when 16#1CCA# => romdata <= X"6C86713C";
    when 16#1CCB# => romdata <= X"43DCDA95";
    when 16#1CCC# => romdata <= X"12B2E717";
    when 16#1CCD# => romdata <= X"3AFC2EF9";
    when 16#1CCE# => romdata <= X"A172C9CF";
    when 16#1CCF# => romdata <= X"DDD3000D";
    when 16#1CD0# => romdata <= X"7A981440";
    when 16#1CD1# => romdata <= X"AD994C39";
    when 16#1CD2# => romdata <= X"DAE6FC0B";
    when 16#1CD3# => romdata <= X"645BA0FD";
    when 16#1CD4# => romdata <= X"49ECAA19";
    when 16#1CD5# => romdata <= X"E572ED0F";
    when 16#1CD6# => romdata <= X"AC748EC8";
    when 16#1CD7# => romdata <= X"37A7D6F2";
    when 16#1CD8# => romdata <= X"8A8D0044";
    when 16#1CD9# => romdata <= X"02F71CA2";
    when 16#1CDA# => romdata <= X"09BB9403";
    when 16#1CDB# => romdata <= X"B21E2983";
    when 16#1CDC# => romdata <= X"6C5FE897";
    when 16#1CDD# => romdata <= X"268DE073";
    when 16#1CDE# => romdata <= X"6E985F96";
    when 16#1CDF# => romdata <= X"31DFDD1A";
    when 16#1CE0# => romdata <= X"C59D5411";
    when 16#1CE1# => romdata <= X"E684BE08";
    when 16#1CE2# => romdata <= X"2F41108E";
    when 16#1CE3# => romdata <= X"33D2B92B";
    when 16#1CE4# => romdata <= X"2D45ED70";
    when 16#1CE5# => romdata <= X"FA52EA2D";
    when 16#1CE6# => romdata <= X"6DE121EB";
    when 16#1CE7# => romdata <= X"9F9C886D";
    when 16#1CE8# => romdata <= X"A479464A";
    when 16#1CE9# => romdata <= X"9DFD9970";
    when 16#1CEA# => romdata <= X"A406491E";
    when 16#1CEB# => romdata <= X"334372D7";
    when 16#1CEC# => romdata <= X"B7893609";
    when 16#1CED# => romdata <= X"5A7459BF";
    when 16#1CEE# => romdata <= X"AFF0E909";
    when 16#1CEF# => romdata <= X"0C2C6B6D";
    when 16#1CF0# => romdata <= X"62624A79";
    when 16#1CF1# => romdata <= X"334F879A";
    when 16#1CF2# => romdata <= X"5C92C685";
    when 16#1CF3# => romdata <= X"B50F75F0";
    when 16#1CF4# => romdata <= X"4BA664EC";
    when 16#1CF5# => romdata <= X"95893FF4";
    when 16#1CF6# => romdata <= X"0D62EEB2";
    when 16#1CF7# => romdata <= X"4DCDD288";
    when 16#1CF8# => romdata <= X"729D0C29";
    when 16#1CF9# => romdata <= X"7DF5ABB8";
    when 16#1CFA# => romdata <= X"3C77FC11";
    when 16#1CFB# => romdata <= X"D0EA3EF1";
    when 16#1CFC# => romdata <= X"8E3BC7C2";
    when 16#1CFD# => romdata <= X"C065CAC5";
    when 16#1CFE# => romdata <= X"1390C610";
    when 16#1CFF# => romdata <= X"B591D240";
    when 16#1D00# => romdata <= X"98CDFCBA";
    when 16#1D01# => romdata <= X"D056240E";
    when 16#1D02# => romdata <= X"180F347C";
    when 16#1D03# => romdata <= X"00912F2D";
    when 16#1D04# => romdata <= X"9ABEBCF5";
    when 16#1D05# => romdata <= X"464D410B";
    when 16#1D06# => romdata <= X"E6A50404";
    when 16#1D07# => romdata <= X"B830F744";
    when 16#1D08# => romdata <= X"D78F7D97";
    when 16#1D09# => romdata <= X"180404FB";
    when 16#1D0A# => romdata <= X"3BCCC228";
    when 16#1D0B# => romdata <= X"8B799181";
    when 16#1D0C# => romdata <= X"0B2562C4";
    when 16#1D0D# => romdata <= X"D509200C";
    when 16#1D0E# => romdata <= X"E1F9C4DF";
    when 16#1D0F# => romdata <= X"6DCA4C60";
    when 16#1D10# => romdata <= X"0D9ED49C";
    when 16#1D11# => romdata <= X"9C145614";
    when 16#1D12# => romdata <= X"1C7B7151";
    when 16#1D13# => romdata <= X"3E728D41";
    when 16#1D14# => romdata <= X"970ACDB6";
    when 16#1D15# => romdata <= X"C15B4A4E";
    when 16#1D16# => romdata <= X"327B9A87";
    when 16#1D17# => romdata <= X"ADA73D1D";
    when 16#1D18# => romdata <= X"46EB0A21";
    when 16#1D19# => romdata <= X"F2F5481C";
    when 16#1D1A# => romdata <= X"3B42931C";
    when 16#1D1B# => romdata <= X"51B780FA";
    when 16#1D1C# => romdata <= X"526C29B9";
    when 16#1D1D# => romdata <= X"8E6B9C71";
    when 16#1D1E# => romdata <= X"4B20049F";
    when 16#1D1F# => romdata <= X"7A05252C";
    when 16#1D20# => romdata <= X"BB84B8E3";
    when 16#1D21# => romdata <= X"6026DB23";
    when 16#1D22# => romdata <= X"79C9632A";
    when 16#1D23# => romdata <= X"0843436E";
    when 16#1D24# => romdata <= X"CB72D15E";
    when 16#1D25# => romdata <= X"A2950ACD";
    when 16#1D26# => romdata <= X"E18DBDC6";
    when 16#1D27# => romdata <= X"DFB01BF0";
    when 16#1D28# => romdata <= X"8F7E191E";
    when 16#1D29# => romdata <= X"C885F11D";
    when 16#1D2A# => romdata <= X"1D8B7BC9";
    when 16#1D2B# => romdata <= X"6E9836B3";
    when 16#1D2C# => romdata <= X"95108F68";
    when 16#1D2D# => romdata <= X"54545082";
    when 16#1D2E# => romdata <= X"A694D597";
    when 16#1D2F# => romdata <= X"4CC36C8A";
    when 16#1D30# => romdata <= X"65834918";
    when 16#1D31# => romdata <= X"6C1BA892";
    when 16#1D32# => romdata <= X"DAA85D3F";
    when 16#1D33# => romdata <= X"156BFBE9";
    when 16#1D34# => romdata <= X"4C73BCD8";
    when 16#1D35# => romdata <= X"15E7652C";
    when 16#1D36# => romdata <= X"38E178AA";
    when 16#1D37# => romdata <= X"F02014F0";
    when 16#1D38# => romdata <= X"E6F23A4E";
    when 16#1D39# => romdata <= X"7EF689EB";
    when 16#1D3A# => romdata <= X"F3ABDCCD";
    when 16#1D3B# => romdata <= X"D40E2DEC";
    when 16#1D3C# => romdata <= X"ED316F07";
    when 16#1D3D# => romdata <= X"E2071692";
    when 16#1D3E# => romdata <= X"7C8F7B20";
    when 16#1D3F# => romdata <= X"3D51D957";
    when 16#1D40# => romdata <= X"EE6EAB06";
    when 16#1D41# => romdata <= X"2B99ACA0";
    when 16#1D42# => romdata <= X"D28E0AB5";
    when 16#1D43# => romdata <= X"0B516CD9";
    when 16#1D44# => romdata <= X"2CBB9BA9";
    when 16#1D45# => romdata <= X"0333E73D";
    when 16#1D46# => romdata <= X"58DE0B4B";
    when 16#1D47# => romdata <= X"633D81EC";
    when 16#1D48# => romdata <= X"93D15EBC";
    when 16#1D49# => romdata <= X"CC813EE6";
    when 16#1D4A# => romdata <= X"3D63BD18";
    when 16#1D4B# => romdata <= X"517F4FE8";
    when 16#1D4C# => romdata <= X"5C374695";
    when 16#1D4D# => romdata <= X"74B8122F";
    when 16#1D4E# => romdata <= X"B9138812";
    when 16#1D4F# => romdata <= X"3E1D5E80";
    when 16#1D50# => romdata <= X"5166FB71";
    when 16#1D51# => romdata <= X"57494F85";
    when 16#1D52# => romdata <= X"59F90A4F";
    when 16#1D53# => romdata <= X"A3DE9E71";
    when 16#1D54# => romdata <= X"DA6FA7CC";
    when 16#1D55# => romdata <= X"C6086E63";
    when 16#1D56# => romdata <= X"8BDD4FD3";
    when 16#1D57# => romdata <= X"E4487506";
    when 16#1D58# => romdata <= X"ACCF84F1";
    when 16#1D59# => romdata <= X"E1678D71";
    when 16#1D5A# => romdata <= X"4B86FAAD";
    when 16#1D5B# => romdata <= X"57A6B76E";
    when 16#1D5C# => romdata <= X"085CFAC3";
    when 16#1D5D# => romdata <= X"0DE469BE";
    when 16#1D5E# => romdata <= X"32E2D203";
    when 16#1D5F# => romdata <= X"C63B43F0";
    when 16#1D60# => romdata <= X"73DD24F4";
    when 16#1D61# => romdata <= X"A1E039B9";
    when 16#1D62# => romdata <= X"41E7A97F";
    when 16#1D63# => romdata <= X"8BB28B51";
    when 16#1D64# => romdata <= X"62174552";
    when 16#1D65# => romdata <= X"68B6EFBB";
    when 16#1D66# => romdata <= X"0E1745C2";
    when 16#1D67# => romdata <= X"3D6D12A8";
    when 16#1D68# => romdata <= X"CD13E5D2";
    when 16#1D69# => romdata <= X"42F562F5";
    when 16#1D6A# => romdata <= X"6FE92496";
    when 16#1D6B# => romdata <= X"342000A7";
    when 16#1D6C# => romdata <= X"31BF3DB0";
    when 16#1D6D# => romdata <= X"A7D31107";
    when 16#1D6E# => romdata <= X"05DFD0D8";
    when 16#1D6F# => romdata <= X"DEFB8566";
    when 16#1D70# => romdata <= X"5B77347C";
    when 16#1D71# => romdata <= X"EFC8629F";
    when 16#1D72# => romdata <= X"3757304F";
    when 16#1D73# => romdata <= X"6129DA98";
    when 16#1D74# => romdata <= X"45F6509F";
    when 16#1D75# => romdata <= X"E3D32DE9";
    when 16#1D76# => romdata <= X"FA86EA4F";
    when 16#1D77# => romdata <= X"A9BF86FF";
    when 16#1D78# => romdata <= X"7CC8E726";
    when 16#1D79# => romdata <= X"C0FA9F93";
    when 16#1D7A# => romdata <= X"F889C467";
    when 16#1D7B# => romdata <= X"642C5E94";
    when 16#1D7C# => romdata <= X"4501BEF8";
    when 16#1D7D# => romdata <= X"ED59793A";
    when 16#1D7E# => romdata <= X"F8804A99";
    when 16#1D7F# => romdata <= X"51B4B880";
    when 16#1D80# => romdata <= X"906F6C5A";
    when 16#1D81# => romdata <= X"1D3BD03A";
    when 16#1D82# => romdata <= X"03802EEF";
    when 16#1D83# => romdata <= X"5937E214";
    when 16#1D84# => romdata <= X"E87B5E2F";
    when 16#1D85# => romdata <= X"0182BA2C";
    when 16#1D86# => romdata <= X"258F44B5";
    when 16#1D87# => romdata <= X"16EC66EA";
    when 16#1D88# => romdata <= X"CB705E06";
    when 16#1D89# => romdata <= X"EA6DFDB5";
    when 16#1D8A# => romdata <= X"6600B846";
    when 16#1D8B# => romdata <= X"3A421DB0";
    when 16#1D8C# => romdata <= X"3A514600";
    when 16#1D8D# => romdata <= X"91D7FE88";
    when 16#1D8E# => romdata <= X"9E6DAE32";
    when 16#1D8F# => romdata <= X"EC19190E";
    when 16#1D90# => romdata <= X"7211F08D";
    when 16#1D91# => romdata <= X"37846CEE";
    when 16#1D92# => romdata <= X"7364B6EC";
    when 16#1D93# => romdata <= X"C07C1740";
    when 16#1D94# => romdata <= X"CE990141";
    when 16#1D95# => romdata <= X"C4DC4CB0";
    when 16#1D96# => romdata <= X"AC9F25CA";
    when 16#1D97# => romdata <= X"FCA6BC91";
    when 16#1D98# => romdata <= X"11102EAB";
    when 16#1D99# => romdata <= X"A250ADFD";
    when 16#1D9A# => romdata <= X"505201FF";
    when 16#1D9B# => romdata <= X"F638B31A";
    when 16#1D9C# => romdata <= X"77CCE7A1";
    when 16#1D9D# => romdata <= X"ECB273F9";
    when 16#1D9E# => romdata <= X"C8ED84EC";
    when 16#1D9F# => romdata <= X"2F403C11";
    when 16#1DA0# => romdata <= X"91596A53";
    when 16#1DA1# => romdata <= X"EAD82342";
    when 16#1DA2# => romdata <= X"1EC47DC5";
    when 16#1DA3# => romdata <= X"E78F3BD1";
    when 16#1DA4# => romdata <= X"339532C9";
    when 16#1DA5# => romdata <= X"7E4EAA02";
    when 16#1DA6# => romdata <= X"4CCC906E";
    when 16#1DA7# => romdata <= X"BFB870C1";
    when 16#1DA8# => romdata <= X"467C3D84";
    when 16#1DA9# => romdata <= X"5A178EB0";
    when 16#1DAA# => romdata <= X"7C11BE8D";
    when 16#1DAB# => romdata <= X"57E4EDEA";
    when 16#1DAC# => romdata <= X"7ADEF162";
    when 16#1DAD# => romdata <= X"923E9521";
    when 16#1DAE# => romdata <= X"451B871D";
    when 16#1DAF# => romdata <= X"F6E357DC";
    when 16#1DB0# => romdata <= X"EEA7F620";
    when 16#1DB1# => romdata <= X"22106F64";
    when 16#1DB2# => romdata <= X"7DD8A230";
    when 16#1DB3# => romdata <= X"74AC10AA";
    when 16#1DB4# => romdata <= X"632C56DC";
    when 16#1DB5# => romdata <= X"32B34A4A";
    when 16#1DB6# => romdata <= X"184FACC6";
    when 16#1DB7# => romdata <= X"4E5D1E8F";
    when 16#1DB8# => romdata <= X"D6926966";
    when 16#1DB9# => romdata <= X"0543EEA2";
    when 16#1DBA# => romdata <= X"FD584117";
    when 16#1DBB# => romdata <= X"A3EBCF62";
    when 16#1DBC# => romdata <= X"68352F02";
    when 16#1DBD# => romdata <= X"12ABCE7C";
    when 16#1DBE# => romdata <= X"D28A93C9";
    when 16#1DBF# => romdata <= X"AF76722F";
    when 16#1DC0# => romdata <= X"B5A71FF9";
    when 16#1DC1# => romdata <= X"E5AC4579";
    when 16#1DC2# => romdata <= X"A2BA32B9";
    when 16#1DC3# => romdata <= X"1818CDCB";
    when 16#1DC4# => romdata <= X"62C77A6A";
    when 16#1DC5# => romdata <= X"8EB1F4C3";
    when 16#1DC6# => romdata <= X"4132EB46";
    when 16#1DC7# => romdata <= X"3812B329";
    when 16#1DC8# => romdata <= X"B6B22108";
    when 16#1DC9# => romdata <= X"AC36E71F";
    when 16#1DCA# => romdata <= X"38338AE3";
    when 16#1DCB# => romdata <= X"A52C6327";
    when 16#1DCC# => romdata <= X"96E45189";
    when 16#1DCD# => romdata <= X"632B73FD";
    when 16#1DCE# => romdata <= X"C0BD37A4";
    when 16#1DCF# => romdata <= X"57204757";
    when 16#1DD0# => romdata <= X"261B7CFC";
    when 16#1DD1# => romdata <= X"01E06BC7";
    when 16#1DD2# => romdata <= X"67A57A5F";
    when 16#1DD3# => romdata <= X"A7CFE437";
    when 16#1DD4# => romdata <= X"94F65398";
    when 16#1DD5# => romdata <= X"A94B4EF0";
    when 16#1DD6# => romdata <= X"9D6DC2A8";
    when 16#1DD7# => romdata <= X"691BD0CB";
    when 16#1DD8# => romdata <= X"018BBE7B";
    when 16#1DD9# => romdata <= X"66E0C37B";
    when 16#1DDA# => romdata <= X"AA472324";
    when 16#1DDB# => romdata <= X"7AF3424B";
    when 16#1DDC# => romdata <= X"DE22614A";
    when 16#1DDD# => romdata <= X"9A581A79";
    when 16#1DDE# => romdata <= X"82E8C232";
    when 16#1DDF# => romdata <= X"3178BD2D";
    when 16#1DE0# => romdata <= X"46E6912A";
    when 16#1DE1# => romdata <= X"2FB2D253";
    when 16#1DE2# => romdata <= X"1819A180";
    when 16#1DE3# => romdata <= X"689D7F2C";
    when 16#1DE4# => romdata <= X"9B5C5AFC";
    when 16#1DE5# => romdata <= X"2DCF1C7F";
    when 16#1DE6# => romdata <= X"AEB1927E";
    when 16#1DE7# => romdata <= X"B79A72EB";
    when 16#1DE8# => romdata <= X"1203BB0F";
    when 16#1DE9# => romdata <= X"F17DAAF2";
    when 16#1DEA# => romdata <= X"7D660221";
    when 16#1DEB# => romdata <= X"95890BBD";
    when 16#1DEC# => romdata <= X"DA786CF1";
    when 16#1DED# => romdata <= X"C36ABFD9";
    when 16#1DEE# => romdata <= X"6BC36FA1";
    when 16#1DEF# => romdata <= X"D2A5A0CC";
    when 16#1DF0# => romdata <= X"3D7EEE1A";
    when 16#1DF1# => romdata <= X"1050CA84";
    when 16#1DF2# => romdata <= X"0209903C";
    when 16#1DF3# => romdata <= X"B9FF429C";
    when 16#1DF4# => romdata <= X"7EE9DF9C";
    when 16#1DF5# => romdata <= X"BC2BAB84";
    when 16#1DF6# => romdata <= X"CF28FAEF";
    when 16#1DF7# => romdata <= X"5BB45AE9";
    when 16#1DF8# => romdata <= X"588970A2";
    when 16#1DF9# => romdata <= X"8B6BD9AD";
    when 16#1DFA# => romdata <= X"F8DF134C";
    when 16#1DFB# => romdata <= X"1FAB0DE2";
    when 16#1DFC# => romdata <= X"74B5C745";
    when 16#1DFD# => romdata <= X"2C4836A5";
    when 16#1DFE# => romdata <= X"73A26A0B";
    when 16#1DFF# => romdata <= X"4C14B740";
    when 16#1E00# => romdata <= X"C6D5046A";
    when 16#1E01# => romdata <= X"5000ECDB";
    when 16#1E02# => romdata <= X"54C872F2";
    when 16#1E03# => romdata <= X"DC494F2D";
    when 16#1E04# => romdata <= X"EB884300";
    when 16#1E05# => romdata <= X"07C9BE8E";
    when 16#1E06# => romdata <= X"C39FFB14";
    when 16#1E07# => romdata <= X"8F00F786";
    when 16#1E08# => romdata <= X"1D827758";
    when 16#1E09# => romdata <= X"9AC839AA";
    when 16#1E0A# => romdata <= X"D30AF7D7";
    when 16#1E0B# => romdata <= X"A2E0F9EE";
    when 16#1E0C# => romdata <= X"8217A39C";
    when 16#1E0D# => romdata <= X"521311E9";
    when 16#1E0E# => romdata <= X"BD59A71B";
    when 16#1E0F# => romdata <= X"C6663A77";
    when 16#1E10# => romdata <= X"38669D6D";
    when 16#1E11# => romdata <= X"3BB28124";
    when 16#1E12# => romdata <= X"A80ABDF9";
    when 16#1E13# => romdata <= X"05DFE2C9";
    when 16#1E14# => romdata <= X"539CCF0C";
    when 16#1E15# => romdata <= X"8FA39EF8";
    when 16#1E16# => romdata <= X"4E9633D6";
    when 16#1E17# => romdata <= X"3BE0C32F";
    when 16#1E18# => romdata <= X"3B2AA9FC";
    when 16#1E19# => romdata <= X"DC18AC38";
    when 16#1E1A# => romdata <= X"C3C00924";
    when 16#1E1B# => romdata <= X"E9D54977";
    when 16#1E1C# => romdata <= X"BDAE6141";
    when 16#1E1D# => romdata <= X"0F997038";
    when 16#1E1E# => romdata <= X"BE066DA6";
    when 16#1E1F# => romdata <= X"C945D825";
    when 16#1E20# => romdata <= X"8B7DD133";
    when 16#1E21# => romdata <= X"EECBA836";
    when 16#1E22# => romdata <= X"A7A6A290";
    when 16#1E23# => romdata <= X"7C431C52";
    when 16#1E24# => romdata <= X"2619D466";
    when 16#1E25# => romdata <= X"430E6ACF";
    when 16#1E26# => romdata <= X"15030F7F";
    when 16#1E27# => romdata <= X"BA4F3D6B";
    when 16#1E28# => romdata <= X"B545CAD8";
    when 16#1E29# => romdata <= X"5678E818";
    when 16#1E2A# => romdata <= X"98D2DE35";
    when 16#1E2B# => romdata <= X"8CFF3951";
    when 16#1E2C# => romdata <= X"C8184066";
    when 16#1E2D# => romdata <= X"B18930DD";
    when 16#1E2E# => romdata <= X"A8678908";
    when 16#1E2F# => romdata <= X"71AF6F41";
    when 16#1E30# => romdata <= X"33B492FC";
    when 16#1E31# => romdata <= X"894DBE4A";
    when 16#1E32# => romdata <= X"A5F1E44B";
    when 16#1E33# => romdata <= X"D361C456";
    when 16#1E34# => romdata <= X"0ABBCD31";
    when 16#1E35# => romdata <= X"01B4AA4E";
    when 16#1E36# => romdata <= X"065FD603";
    when 16#1E37# => romdata <= X"08795DDA";
    when 16#1E38# => romdata <= X"EBADBB60";
    when 16#1E39# => romdata <= X"4A3D5877";
    when 16#1E3A# => romdata <= X"6006CD07";
    when 16#1E3B# => romdata <= X"4389AF49";
    when 16#1E3C# => romdata <= X"A0EF0958";
    when 16#1E3D# => romdata <= X"6410015C";
    when 16#1E3E# => romdata <= X"7DE4FEFE";
    when 16#1E3F# => romdata <= X"EBEA6262";
    when 16#1E40# => romdata <= X"B23571B9";
    when 16#1E41# => romdata <= X"3BEE15CD";
    when 16#1E42# => romdata <= X"A2BBA60B";
    when 16#1E43# => romdata <= X"6CC72A7D";
    when 16#1E44# => romdata <= X"C9C80C81";
    when 16#1E45# => romdata <= X"C9A25FE3";
    when 16#1E46# => romdata <= X"D149C7A8";
    when 16#1E47# => romdata <= X"BB2F704B";
    when 16#1E48# => romdata <= X"E11177F9";
    when 16#1E49# => romdata <= X"2E2CEF0B";
    when 16#1E4A# => romdata <= X"BD12C076";
    when 16#1E4B# => romdata <= X"6D691CCF";
    when 16#1E4C# => romdata <= X"093D456A";
    when 16#1E4D# => romdata <= X"FEA411A8";
    when 16#1E4E# => romdata <= X"FE5F1C1A";
    when 16#1E4F# => romdata <= X"44F31017";
    when 16#1E50# => romdata <= X"760F0D0C";
    when 16#1E51# => romdata <= X"C3B271FB";
    when 16#1E52# => romdata <= X"15F56D9F";
    when 16#1E53# => romdata <= X"51A594C3";
    when 16#1E54# => romdata <= X"4FDFF8F8";
    when 16#1E55# => romdata <= X"ADC91584";
    when 16#1E56# => romdata <= X"ED8D7E1B";
    when 16#1E57# => romdata <= X"6DAB27B2";
    when 16#1E58# => romdata <= X"BE1BBDC4";
    when 16#1E59# => romdata <= X"486FB1C8";
    when 16#1E5A# => romdata <= X"22F23704";
    when 16#1E5B# => romdata <= X"BB2EF4B5";
    when 16#1E5C# => romdata <= X"21E02E42";
    when 16#1E5D# => romdata <= X"FDCABF69";
    when 16#1E5E# => romdata <= X"588B0B9D";
    when 16#1E5F# => romdata <= X"92AAA731";
    when 16#1E60# => romdata <= X"16D26E8E";
    when 16#1E61# => romdata <= X"9E48DE94";
    when 16#1E62# => romdata <= X"F6267414";
    when 16#1E63# => romdata <= X"AC845467";
    when 16#1E64# => romdata <= X"597B4C1F";
    when 16#1E65# => romdata <= X"2A9A8E1E";
    when 16#1E66# => romdata <= X"82C0A1C0";
    when 16#1E67# => romdata <= X"5955022C";
    when 16#1E68# => romdata <= X"DF873860";
    when 16#1E69# => romdata <= X"98EAFC5B";
    when 16#1E6A# => romdata <= X"F1A04071";
    when 16#1E6B# => romdata <= X"6A89BE53";
    when 16#1E6C# => romdata <= X"A36B1433";
    when 16#1E6D# => romdata <= X"76927028";
    when 16#1E6E# => romdata <= X"A561BBC0";
    when 16#1E6F# => romdata <= X"7AFAF424";
    when 16#1E70# => romdata <= X"94DF5BC0";
    when 16#1E71# => romdata <= X"D95170D8";
    when 16#1E72# => romdata <= X"53DCCCCB";
    when 16#1E73# => romdata <= X"22FD36B7";
    when 16#1E74# => romdata <= X"947712EB";
    when 16#1E75# => romdata <= X"369077D0";
    when 16#1E76# => romdata <= X"2BF85B0A";
    when 16#1E77# => romdata <= X"4F57757E";
    when 16#1E78# => romdata <= X"D80B247E";
    when 16#1E79# => romdata <= X"521AC640";
    when 16#1E7A# => romdata <= X"D1B1CE30";
    when 16#1E7B# => romdata <= X"F93DEBBE";
    when 16#1E7C# => romdata <= X"2389D364";
    when 16#1E7D# => romdata <= X"A8B7971A";
    when 16#1E7E# => romdata <= X"51AFA4F5";
    when 16#1E7F# => romdata <= X"57A8E120";
    when 16#1E80# => romdata <= X"FDCF36E6";
    when 16#1E81# => romdata <= X"C842D2AB";
    when 16#1E82# => romdata <= X"CCE9D878";
    when 16#1E83# => romdata <= X"3D0D7A7E";
    when 16#1E84# => romdata <= X"B74992EA";
    when 16#1E85# => romdata <= X"CEEF6C61";
    when 16#1E86# => romdata <= X"8AC7DED4";
    when 16#1E87# => romdata <= X"E457B1A7";
    when 16#1E88# => romdata <= X"08BE2C82";
    when 16#1E89# => romdata <= X"B28A9563";
    when 16#1E8A# => romdata <= X"F4A088FF";
    when 16#1E8B# => romdata <= X"7DB146B1";
    when 16#1E8C# => romdata <= X"6B47A900";
    when 16#1E8D# => romdata <= X"DF49A4F3";
    when 16#1E8E# => romdata <= X"FA8EDAAF";
    when 16#1E8F# => romdata <= X"CA09F408";
    when 16#1E90# => romdata <= X"B025D04E";
    when 16#1E91# => romdata <= X"B673E105";
    when 16#1E92# => romdata <= X"E0F55959";
    when 16#1E93# => romdata <= X"B7951CF0";
    when 16#1E94# => romdata <= X"E999CDF6";
    when 16#1E95# => romdata <= X"8EA9B323";
    when 16#1E96# => romdata <= X"33DBFE05";
    when 16#1E97# => romdata <= X"16D27211";
    when 16#1E98# => romdata <= X"1CBBD993";
    when 16#1E99# => romdata <= X"3CA8AD8A";
    when 16#1E9A# => romdata <= X"A6025E5F";
    when 16#1E9B# => romdata <= X"9A062D83";
    when 16#1E9C# => romdata <= X"05344CAF";
    when 16#1E9D# => romdata <= X"C3CA391B";
    when 16#1E9E# => romdata <= X"D8DEBDC5";
    when 16#1E9F# => romdata <= X"8F7FDBC0";
    when 16#1EA0# => romdata <= X"41B34990";
    when 16#1EA1# => romdata <= X"0E397609";
    when 16#1EA2# => romdata <= X"C71E4EA3";
    when 16#1EA3# => romdata <= X"A9D8407C";
    when 16#1EA4# => romdata <= X"63E8A6BB";
    when 16#1EA5# => romdata <= X"EEAEFC92";
    when 16#1EA6# => romdata <= X"E9C93914";
    when 16#1EA7# => romdata <= X"7920E48E";
    when 16#1EA8# => romdata <= X"35DAC6D1";
    when 16#1EA9# => romdata <= X"23DA46E4";
    when 16#1EAA# => romdata <= X"F0838FD7";
    when 16#1EAB# => romdata <= X"32E43FE4";
    when 16#1EAC# => romdata <= X"EEF6BD68";
    when 16#1EAD# => romdata <= X"D5AF0C9B";
    when 16#1EAE# => romdata <= X"A3A0CB28";
    when 16#1EAF# => romdata <= X"233743B2";
    when 16#1EB0# => romdata <= X"91D4E100";
    when 16#1EB1# => romdata <= X"54F695DC";
    when 16#1EB2# => romdata <= X"10A847E6";
    when 16#1EB3# => romdata <= X"61F39C4C";
    when 16#1EB4# => romdata <= X"133289B0";
    when 16#1EB5# => romdata <= X"7ACA8B54";
    when 16#1EB6# => romdata <= X"4EE3E2EC";
    when 16#1EB7# => romdata <= X"288CB18C";
    when 16#1EB8# => romdata <= X"40CD9A8E";
    when 16#1EB9# => romdata <= X"48A93378";
    when 16#1EBA# => romdata <= X"FD50E077";
    when 16#1EBB# => romdata <= X"EFBC2199";
    when 16#1EBC# => romdata <= X"6424B539";
    when 16#1EBD# => romdata <= X"A397B3D2";
    when 16#1EBE# => romdata <= X"A6C7DE58";
    when 16#1EBF# => romdata <= X"112CF55E";
    when 16#1EC0# => romdata <= X"82E8FF10";
    when 16#1EC1# => romdata <= X"F75571A1";
    when 16#1EC2# => romdata <= X"5DC248E6";
    when 16#1EC3# => romdata <= X"B77CBB91";
    when 16#1EC4# => romdata <= X"D8BF2D53";
    when 16#1EC5# => romdata <= X"E5C4E9A8";
    when 16#1EC6# => romdata <= X"5C7EB8FB";
    when 16#1EC7# => romdata <= X"690F74BE";
    when 16#1EC8# => romdata <= X"029CE1B5";
    when 16#1EC9# => romdata <= X"69EFACFC";
    when 16#1ECA# => romdata <= X"16872C50";
    when 16#1ECB# => romdata <= X"08820FC6";
    when 16#1ECC# => romdata <= X"A7D12AB4";
    when 16#1ECD# => romdata <= X"3E08B4AF";
    when 16#1ECE# => romdata <= X"F57DE6B4";
    when 16#1ECF# => romdata <= X"3B613DF8";
    when 16#1ED0# => romdata <= X"480ACA55";
    when 16#1ED1# => romdata <= X"6E29D792";
    when 16#1ED2# => romdata <= X"C6C81CB1";
    when 16#1ED3# => romdata <= X"CB54A672";
    when 16#1ED4# => romdata <= X"45C571A0";
    when 16#1ED5# => romdata <= X"4965267B";
    when 16#1ED6# => romdata <= X"A0F9CD3F";
    when 16#1ED7# => romdata <= X"A0950B9A";
    when 16#1ED8# => romdata <= X"5B393B4A";
    when 16#1ED9# => romdata <= X"230A41E4";
    when 16#1EDA# => romdata <= X"55267CD3";
    when 16#1EDB# => romdata <= X"96F42285";
    when 16#1EDC# => romdata <= X"F0E49C5A";
    when 16#1EDD# => romdata <= X"FA0B53EC";
    when 16#1EDE# => romdata <= X"7B60C1C3";
    when 16#1EDF# => romdata <= X"17EDA3FA";
    when 16#1EE0# => romdata <= X"E4B1713A";
    when 16#1EE1# => romdata <= X"80D4EBAD";
    when 16#1EE2# => romdata <= X"32FC685C";
    when 16#1EE3# => romdata <= X"13649C48";
    when 16#1EE4# => romdata <= X"06D6FD88";
    when 16#1EE5# => romdata <= X"7A24A4F7";
    when 16#1EE6# => romdata <= X"AE801405";
    when 16#1EE7# => romdata <= X"EF28F058";
    when 16#1EE8# => romdata <= X"B37112A6";
    when 16#1EE9# => romdata <= X"80F9E9AD";
    when 16#1EEA# => romdata <= X"0456314E";
    when 16#1EEB# => romdata <= X"9F490393";
    when 16#1EEC# => romdata <= X"CA257757";
    when 16#1EED# => romdata <= X"97E4CCF9";
    when 16#1EEE# => romdata <= X"184FF0C6";
    when 16#1EEF# => romdata <= X"A237AFFA";
    when 16#1EF0# => romdata <= X"8DE1B84C";
    when 16#1EF1# => romdata <= X"420A6183";
    when 16#1EF2# => romdata <= X"B1D49D6F";
    when 16#1EF3# => romdata <= X"2AC1E673";
    when 16#1EF4# => romdata <= X"E7FDE161";
    when 16#1EF5# => romdata <= X"A8159DCE";
    when 16#1EF6# => romdata <= X"B00D85F0";
    when 16#1EF7# => romdata <= X"32EE76E3";
    when 16#1EF8# => romdata <= X"931C459C";
    when 16#1EF9# => romdata <= X"E935DFE4";
    when 16#1EFA# => romdata <= X"AD6C6110";
    when 16#1EFB# => romdata <= X"591EE584";
    when 16#1EFC# => romdata <= X"96B82A16";
    when 16#1EFD# => romdata <= X"630E8232";
    when 16#1EFE# => romdata <= X"0B951088";
    when 16#1EFF# => romdata <= X"0BE4E720";
    when 16#1F00# => romdata <= X"94964FC9";
    when 16#1F01# => romdata <= X"F66389FE";
    when 16#1F02# => romdata <= X"3880283C";
    when 16#1F03# => romdata <= X"4250E6E1";
    when 16#1F04# => romdata <= X"9F195DFE";
    when 16#1F05# => romdata <= X"BD2104FC";
    when 16#1F06# => romdata <= X"0959E084";
    when 16#1F07# => romdata <= X"308BC9CF";
    when 16#1F08# => romdata <= X"DC6E5ED1";
    when 16#1F09# => romdata <= X"C4B48B4E";
    when 16#1F0A# => romdata <= X"CAEB4FDE";
    when 16#1F0B# => romdata <= X"5F215FBE";
    when 16#1F0C# => romdata <= X"D85A6CD4";
    when 16#1F0D# => romdata <= X"D1C1466E";
    when 16#1F0E# => romdata <= X"68A4CF21";
    when 16#1F0F# => romdata <= X"AEF29F77";
    when 16#1F10# => romdata <= X"933549A3";
    when 16#1F11# => romdata <= X"A6FF7ACD";
    when 16#1F12# => romdata <= X"8AB6E6C6";
    when 16#1F13# => romdata <= X"89F1E8DF";
    when 16#1F14# => romdata <= X"0AD8AB28";
    when 16#1F15# => romdata <= X"9D5C3302";
    when 16#1F16# => romdata <= X"3DF90B21";
    when 16#1F17# => romdata <= X"A26320CE";
    when 16#1F18# => romdata <= X"8C1CEB2C";
    when 16#1F19# => romdata <= X"099FC1DB";
    when 16#1F1A# => romdata <= X"58737665";
    when 16#1F1B# => romdata <= X"855DCD20";
    when 16#1F1C# => romdata <= X"D587E176";
    when 16#1F1D# => romdata <= X"483E33EF";
    when 16#1F1E# => romdata <= X"14C80AA4";
    when 16#1F1F# => romdata <= X"760F751E";
    when 16#1F20# => romdata <= X"E5B28460";
    when 16#1F21# => romdata <= X"811E5110";
    when 16#1F22# => romdata <= X"FEC3D689";
    when 16#1F23# => romdata <= X"AE2A6E91";
    when 16#1F24# => romdata <= X"D0A3F1E2";
    when 16#1F25# => romdata <= X"2623E885";
    when 16#1F26# => romdata <= X"71F4DAC8";
    when 16#1F27# => romdata <= X"95AA428D";
    when 16#1F28# => romdata <= X"42634EC1";
    when 16#1F29# => romdata <= X"42E56D0D";
    when 16#1F2A# => romdata <= X"57CE68D7";
    when 16#1F2B# => romdata <= X"949BE13A";
    when 16#1F2C# => romdata <= X"F234229E";
    when 16#1F2D# => romdata <= X"546E9D66";
    when 16#1F2E# => romdata <= X"D5C58E51";
    when 16#1F2F# => romdata <= X"0BF3EAC7";
    when 16#1F30# => romdata <= X"B73309BE";
    when 16#1F31# => romdata <= X"16DCE6E2";
    when 16#1F32# => romdata <= X"280AA802";
    when 16#1F33# => romdata <= X"47D9EDED";
    when 16#1F34# => romdata <= X"D20E0629";
    when 16#1F35# => romdata <= X"5C9876B4";
    when 16#1F36# => romdata <= X"12B786CF";
    when 16#1F37# => romdata <= X"7E5F1073";
    when 16#1F38# => romdata <= X"79215813";
    when 16#1F39# => romdata <= X"1AFA002F";
    when 16#1F3A# => romdata <= X"E7750A17";
    when 16#1F3B# => romdata <= X"015A9C25";
    when 16#1F3C# => romdata <= X"80646A9A";
    when 16#1F3D# => romdata <= X"0D2A3F02";
    when 16#1F3E# => romdata <= X"43AF1AB4";
    when 16#1F3F# => romdata <= X"FEFB3D02";
    when 16#1F40# => romdata <= X"8504553A";
    when 16#1F41# => romdata <= X"F9C5C34D";
    when 16#1F42# => romdata <= X"1A4A2FE3";
    when 16#1F43# => romdata <= X"B8DD8BF8";
    when 16#1F44# => romdata <= X"CEADA82A";
    when 16#1F45# => romdata <= X"E63C319B";
    when 16#1F46# => romdata <= X"D7981D97";
    when 16#1F47# => romdata <= X"155AA2F1";
    when 16#1F48# => romdata <= X"05D724A8";
    when 16#1F49# => romdata <= X"C09310D5";
    when 16#1F4A# => romdata <= X"C3168770";
    when 16#1F4B# => romdata <= X"62152419";
    when 16#1F4C# => romdata <= X"A006ABF5";
    when 16#1F4D# => romdata <= X"6AADED74";
    when 16#1F4E# => romdata <= X"DF0DF325";
    when 16#1F4F# => romdata <= X"D666C31D";
    when 16#1F50# => romdata <= X"F51F194C";
    when 16#1F51# => romdata <= X"FEB331E7";
    when 16#1F52# => romdata <= X"DAF00410";
    when 16#1F53# => romdata <= X"372999D2";
    when 16#1F54# => romdata <= X"D05B023B";
    when 16#1F55# => romdata <= X"2C3067E6";
    when 16#1F56# => romdata <= X"CE4A472F";
    when 16#1F57# => romdata <= X"ED3B8BE1";
    when 16#1F58# => romdata <= X"C15C24DF";
    when 16#1F59# => romdata <= X"BF4956A5";
    when 16#1F5A# => romdata <= X"B670FFCF";
    when 16#1F5B# => romdata <= X"128E5A23";
    when 16#1F5C# => romdata <= X"039764BE";
    when 16#1F5D# => romdata <= X"39CBE556";
    when 16#1F5E# => romdata <= X"36B83674";
    when 16#1F5F# => romdata <= X"060B3CCF";
    when 16#1F60# => romdata <= X"5EF9A7B7";
    when 16#1F61# => romdata <= X"EAB0813A";
    when 16#1F62# => romdata <= X"DEE82E27";
    when 16#1F63# => romdata <= X"1C422FB7";
    when 16#1F64# => romdata <= X"8A982000";
    when 16#1F65# => romdata <= X"7753B1E6";
    when 16#1F66# => romdata <= X"2BF4CCC0";
    when 16#1F67# => romdata <= X"74F7796D";
    when 16#1F68# => romdata <= X"5B2008FE";
    when 16#1F69# => romdata <= X"6542DC0C";
    when 16#1F6A# => romdata <= X"77ECA381";
    when 16#1F6B# => romdata <= X"0120ABE9";
    when 16#1F6C# => romdata <= X"F90BE593";
    when 16#1F6D# => romdata <= X"4E8EAE36";
    when 16#1F6E# => romdata <= X"5D02B3D2";
    when 16#1F6F# => romdata <= X"DF4EA4A8";
    when 16#1F70# => romdata <= X"27E03326";
    when 16#1F71# => romdata <= X"3B113EEE";
    when 16#1F72# => romdata <= X"5823DD39";
    when 16#1F73# => romdata <= X"12FB31E3";
    when 16#1F74# => romdata <= X"C4B46B27";
    when 16#1F75# => romdata <= X"4D7115F3";
    when 16#1F76# => romdata <= X"4CDA793D";
    when 16#1F77# => romdata <= X"B6AD2CD8";
    when 16#1F78# => romdata <= X"BCAF4B13";
    when 16#1F79# => romdata <= X"B832AB60";
    when 16#1F7A# => romdata <= X"5BE42B28";
    when 16#1F7B# => romdata <= X"77EE2E66";
    when 16#1F7C# => romdata <= X"B411668E";
    when 16#1F7D# => romdata <= X"A29A7DBA";
    when 16#1F7E# => romdata <= X"5BD969B9";
    when 16#1F7F# => romdata <= X"F1526380";
    when 16#1F80# => romdata <= X"9B8071D9";
    when 16#1F81# => romdata <= X"6E7D361B";
    when 16#1F82# => romdata <= X"2462CA93";
    when 16#1F83# => romdata <= X"748DE4D3";
    when 16#1F84# => romdata <= X"1746972D";
    when 16#1F85# => romdata <= X"AE582AD4";
    when 16#1F86# => romdata <= X"F70A188C";
    when 16#1F87# => romdata <= X"B40C2E6E";
    when 16#1F88# => romdata <= X"418288B6";
    when 16#1F89# => romdata <= X"A713ED4B";
    when 16#1F8A# => romdata <= X"647013B3";
    when 16#1F8B# => romdata <= X"EC31C9EA";
    when 16#1F8C# => romdata <= X"6217DE55";
    when 16#1F8D# => romdata <= X"D016A197";
    when 16#1F8E# => romdata <= X"7A0B2852";
    when 16#1F8F# => romdata <= X"24129CDC";
    when 16#1F90# => romdata <= X"59A9E54F";
    when 16#1F91# => romdata <= X"3E509425";
    when 16#1F92# => romdata <= X"8F11C0C9";
    when 16#1F93# => romdata <= X"95F60785";
    when 16#1F94# => romdata <= X"614E5607";
    when 16#1F95# => romdata <= X"64312CD8";
    when 16#1F96# => romdata <= X"6C6969B3";
    when 16#1F97# => romdata <= X"274236EE";
    when 16#1F98# => romdata <= X"602EFAE3";
    when 16#1F99# => romdata <= X"92C015E4";
    when 16#1F9A# => romdata <= X"C3972D6F";
    when 16#1F9B# => romdata <= X"A2A47AB4";
    when 16#1F9C# => romdata <= X"8D5C5F68";
    when 16#1F9D# => romdata <= X"36AFA54F";
    when 16#1F9E# => romdata <= X"28CCC03B";
    when 16#1F9F# => romdata <= X"B4DAA0A1";
    when 16#1FA0# => romdata <= X"DC0DCA3F";
    when 16#1FA1# => romdata <= X"D3F2B15F";
    when 16#1FA2# => romdata <= X"B2ADD907";
    when 16#1FA3# => romdata <= X"D3BF7719";
    when 16#1FA4# => romdata <= X"D1D9A828";
    when 16#1FA5# => romdata <= X"4A47C30F";
    when 16#1FA6# => romdata <= X"32712A8C";
    when 16#1FA7# => romdata <= X"D440148B";
    when 16#1FA8# => romdata <= X"8DFDB851";
    when 16#1FA9# => romdata <= X"FFD25ECA";
    when 16#1FAA# => romdata <= X"2864150B";
    when 16#1FAB# => romdata <= X"832F8B5D";
    when 16#1FAC# => romdata <= X"C3A7C701";
    when 16#1FAD# => romdata <= X"371785A6";
    when 16#1FAE# => romdata <= X"6285601E";
    when 16#1FAF# => romdata <= X"96D285FF";
    when 16#1FB0# => romdata <= X"88947804";
    when 16#1FB1# => romdata <= X"AA4D8866";
    when 16#1FB2# => romdata <= X"5B3E1576";
    when 16#1FB3# => romdata <= X"0CDE327F";
    when 16#1FB4# => romdata <= X"BD213930";
    when 16#1FB5# => romdata <= X"42BAF62F";
    when 16#1FB6# => romdata <= X"DCE6EC41";
    when 16#1FB7# => romdata <= X"955E877E";
    when 16#1FB8# => romdata <= X"CAC331D5";
    when 16#1FB9# => romdata <= X"94ED4054";
    when 16#1FBA# => romdata <= X"7AFED34D";
    when 16#1FBB# => romdata <= X"410714CE";
    when 16#1FBC# => romdata <= X"57FCB4F0";
    when 16#1FBD# => romdata <= X"1C882651";
    when 16#1FBE# => romdata <= X"9ACB85F4";
    when 16#1FBF# => romdata <= X"47306C86";
    when 16#1FC0# => romdata <= X"BD1BA818";
    when 16#1FC1# => romdata <= X"9E0621DD";
    when 16#1FC2# => romdata <= X"09451E8F";
    when 16#1FC3# => romdata <= X"341AE47E";
    when 16#1FC4# => romdata <= X"7FCF1FD2";
    when 16#1FC5# => romdata <= X"DE2AF78E";
    when 16#1FC6# => romdata <= X"0AFA27A4";
    when 16#1FC7# => romdata <= X"B6DD51A0";
    when 16#1FC8# => romdata <= X"710FC1FC";
    when 16#1FC9# => romdata <= X"4A599823";
    when 16#1FCA# => romdata <= X"4EDAA1D4";
    when 16#1FCB# => romdata <= X"CF0786B7";
    when 16#1FCC# => romdata <= X"79F637EE";
    when 16#1FCD# => romdata <= X"1A720587";
    when 16#1FCE# => romdata <= X"74C1B4BF";
    when 16#1FCF# => romdata <= X"5E125DEB";
    when 16#1FD0# => romdata <= X"B4230645";
    when 16#1FD1# => romdata <= X"ECF87E3C";
    when 16#1FD2# => romdata <= X"6FDC91E1";
    when 16#1FD3# => romdata <= X"D14397FA";
    when 16#1FD4# => romdata <= X"72686784";
    when 16#1FD5# => romdata <= X"815D9654";
    when 16#1FD6# => romdata <= X"839AE8FA";
    when 16#1FD7# => romdata <= X"43864709";
    when 16#1FD8# => romdata <= X"EE0F4A33";
    when 16#1FD9# => romdata <= X"6E3C399C";
    when 16#1FDA# => romdata <= X"A20B2E65";
    when 16#1FDB# => romdata <= X"2E2AB177";
    when 16#1FDC# => romdata <= X"19F9253F";
    when 16#1FDD# => romdata <= X"772EB7A9";
    when 16#1FDE# => romdata <= X"E8838FED";
    when 16#1FDF# => romdata <= X"4EBCD0F8";
    when 16#1FE0# => romdata <= X"CD977583";
    when 16#1FE1# => romdata <= X"BDCEEBBD";
    when 16#1FE2# => romdata <= X"925676F5";
    when 16#1FE3# => romdata <= X"6AAB0C36";
    when 16#1FE4# => romdata <= X"F3DD915F";
    when 16#1FE5# => romdata <= X"6691A30D";
    when 16#1FE6# => romdata <= X"60D52321";
    when 16#1FE7# => romdata <= X"6FB233CB";
    when 16#1FE8# => romdata <= X"BEDE7FDF";
    when 16#1FE9# => romdata <= X"BA827450";
    when 16#1FEA# => romdata <= X"E595AB51";
    when 16#1FEB# => romdata <= X"237F9E77";
    when 16#1FEC# => romdata <= X"058E40F8";
    when 16#1FED# => romdata <= X"62D3A5A9";
    when 16#1FEE# => romdata <= X"6E4AA3DA";
    when 16#1FEF# => romdata <= X"74503812";
    when 16#1FF0# => romdata <= X"EDEFA501";
    when 16#1FF1# => romdata <= X"E526DB6B";
    when 16#1FF2# => romdata <= X"4C642222";
    when 16#1FF3# => romdata <= X"D7F33B06";
    when 16#1FF4# => romdata <= X"D9CD0023";
    when 16#1FF5# => romdata <= X"471DF573";
    when 16#1FF6# => romdata <= X"0CF8E2BE";
    when 16#1FF7# => romdata <= X"E834D108";
    when 16#1FF8# => romdata <= X"A25729C1";
    when 16#1FF9# => romdata <= X"C1484C20";
    when 16#1FFA# => romdata <= X"7ECEB0E4";
    when 16#1FFB# => romdata <= X"598965EA";
    when 16#1FFC# => romdata <= X"B5216D4E";
    when 16#1FFD# => romdata <= X"7C30577A";
    when 16#1FFE# => romdata <= X"89FB8BEC";
    when 16#1FFF# => romdata <= X"0B118F40";
    when others => romdata <= (others => '0');
    end case;
  end process;
end;
